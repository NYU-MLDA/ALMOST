//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT8), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT9), .ZN(new_n229_));
  AOI211_X1 g028(.A(new_n229_), .B(new_n219_), .C1(KEYINPUT9), .C2(new_n213_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n221_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n212_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT67), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n210_), .B(KEYINPUT65), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n236_), .A2(new_n237_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT66), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n203_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT12), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n210_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(KEYINPUT12), .A3(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n243_), .A2(new_n202_), .A3(new_n245_), .A4(new_n239_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G120gat), .B(G148gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(G176gat), .B(G204gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n241_), .A2(new_n246_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n256_));
  NAND2_X1  g055(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI22_X1  g057(.A1(new_n254_), .A2(new_n255_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n255_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n253_), .A3(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263_));
  INV_X1    g062(.A(G1gat), .ZN(new_n264_));
  INV_X1    g063(.A(G8gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n263_), .B1(new_n266_), .B2(KEYINPUT72), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(KEYINPUT72), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G1gat), .B(G8gat), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(G231gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(new_n210_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT17), .ZN(new_n277_));
  XOR2_X1   g076(.A(G127gat), .B(G155gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT16), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G183gat), .B(G211gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n276_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(new_n274_), .B2(new_n244_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n212_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n235_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n281_), .B(KEYINPUT17), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G29gat), .B(G36gat), .Z(new_n290_));
  XOR2_X1   g089(.A(G43gat), .B(G50gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G232gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT34), .ZN(new_n295_));
  OAI22_X1  g094(.A1(new_n232_), .A2(new_n293_), .B1(KEYINPUT35), .B2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n292_), .B(KEYINPUT15), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n232_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(KEYINPUT35), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G190gat), .B(G218gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT70), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT36), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n300_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n301_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n305_), .A2(KEYINPUT36), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n306_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT71), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n307_), .B2(new_n301_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT37), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n301_), .A2(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n311_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT37), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n308_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n262_), .A2(new_n289_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n320_), .B(KEYINPUT73), .Z(new_n321_));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n325_), .A2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n324_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n327_), .A3(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT31), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n350_));
  NOR2_X1   g149(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n337_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(KEYINPUT23), .B2(new_n337_), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n354_), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G190gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT25), .B1(new_n354_), .B2(KEYINPUT76), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n353_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n349_), .A2(new_n364_), .A3(KEYINPUT30), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT30), .B1(new_n349_), .B2(new_n364_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT30), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n353_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n342_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n347_), .B1(new_n370_), .B2(new_n341_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n349_), .A2(new_n364_), .A3(KEYINPUT30), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n367_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G15gat), .B(G43gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(G71gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G99gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n383_), .B(G99gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n379_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n372_), .A2(new_n374_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(KEYINPUT80), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n335_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n389_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n367_), .B2(new_n375_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n396_), .A2(new_n392_), .A3(new_n334_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n322_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n393_), .A3(new_n335_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n334_), .B1(new_n396_), .B2(new_n392_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT82), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT21), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G211gat), .B(G218gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT85), .ZN(new_n407_));
  INV_X1    g206(.A(G204gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n410_));
  NAND2_X1  g209(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(G197gat), .A4(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G197gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT84), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G197gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n416_), .A3(G204gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n409_), .A2(G197gat), .A3(new_n411_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT86), .ZN(new_n420_));
  AOI211_X1 g219(.A(new_n405_), .B(new_n406_), .C1(new_n418_), .C2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(new_n405_), .A3(new_n417_), .A4(new_n412_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n418_), .A2(KEYINPUT87), .A3(new_n405_), .A4(new_n420_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(new_n416_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n409_), .A2(new_n411_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n427_), .A2(new_n408_), .B1(new_n428_), .B2(new_n413_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n406_), .B1(new_n429_), .B2(new_n405_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n421_), .B1(new_n426_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433_));
  NAND3_X1  g232(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT1), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT1), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n434_), .ZN(new_n442_));
  INV_X1    g241(.A(G155gat), .ZN(new_n443_));
  INV_X1    g242(.A(G162gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G141gat), .A2(G148gat), .ZN(new_n447_));
  INV_X1    g246(.A(G141gat), .ZN(new_n448_));
  INV_X1    g247(.A(G148gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n447_), .B(KEYINPUT2), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n450_), .A2(KEYINPUT3), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(KEYINPUT3), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n440_), .A2(new_n434_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n433_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n404_), .B1(new_n432_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n458_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n430_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n460_), .B(new_n403_), .C1(new_n461_), .C2(new_n421_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G78gat), .B(G106gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466_));
  INV_X1    g265(.A(new_n464_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n462_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n451_), .A2(new_n457_), .A3(new_n433_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT28), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT28), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n451_), .A2(new_n457_), .A3(new_n472_), .A4(new_n433_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G22gat), .B(G50gat), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n459_), .A2(KEYINPUT88), .A3(new_n462_), .A4(new_n467_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n469_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n468_), .A2(new_n477_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n467_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n465_), .A2(KEYINPUT89), .A3(new_n468_), .A4(new_n477_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n402_), .A2(new_n480_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G8gat), .B(G36gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G64gat), .B(G92gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n492_), .A2(KEYINPUT32), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n349_), .A2(new_n364_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n461_), .A2(new_n494_), .A3(new_n421_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT91), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n426_), .A2(new_n431_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n421_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT20), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n498_), .A2(new_n500_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT25), .B(G183gat), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n356_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n363_), .A3(new_n370_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT22), .B(G169gat), .Z(new_n513_));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT22), .B(G169gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT93), .ZN(new_n517_));
  AOI21_X1  g316(.A(G176gat), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n362_), .B(KEYINPUT92), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n521_), .B2(new_n340_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n512_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n508_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n497_), .A2(new_n503_), .A3(new_n507_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n508_), .A2(KEYINPUT94), .A3(new_n494_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n432_), .B2(new_n499_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n523_), .A2(KEYINPUT97), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT97), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n512_), .B(new_n532_), .C1(new_n518_), .C2(new_n522_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n496_), .B1(new_n534_), .B2(new_n432_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n507_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n493_), .B1(new_n526_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n451_), .A2(new_n457_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n333_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n451_), .A2(new_n332_), .A3(new_n330_), .A4(new_n457_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(KEYINPUT4), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n333_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n538_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G1gat), .B(G29gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G85gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT0), .B(G57gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n538_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n545_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n497_), .A2(new_n503_), .A3(new_n524_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n523_), .ZN(new_n556_));
  AOI211_X1 g355(.A(new_n496_), .B(new_n506_), .C1(new_n432_), .C2(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n555_), .A2(new_n506_), .B1(new_n530_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n493_), .B(KEYINPUT96), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n537_), .B(new_n554_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT33), .B(new_n549_), .C1(new_n545_), .C2(new_n551_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n542_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n549_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n540_), .A2(new_n550_), .A3(new_n541_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n563_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n496_), .B1(new_n432_), .B2(new_n499_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n570_), .A2(new_n502_), .B1(new_n508_), .B2(new_n523_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n507_), .B1(new_n571_), .B2(new_n497_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n530_), .A2(new_n557_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n491_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n555_), .A2(new_n506_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n530_), .A2(new_n557_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n492_), .A3(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n486_), .B1(new_n561_), .B2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT27), .B1(new_n574_), .B2(new_n577_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n531_), .A2(new_n533_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT20), .B1(new_n582_), .B2(new_n508_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n529_), .B2(new_n527_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n525_), .B1(new_n584_), .B2(new_n507_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n581_), .B1(new_n585_), .B2(new_n491_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n577_), .A2(KEYINPUT27), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n581_), .A3(new_n491_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n580_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n484_), .A2(new_n485_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n478_), .A2(new_n479_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n483_), .A2(KEYINPUT88), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n593_), .B2(new_n468_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n402_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n394_), .A2(new_n397_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n480_), .A2(new_n596_), .A3(new_n484_), .A4(new_n485_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n554_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n579_), .B1(new_n590_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT75), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n272_), .A2(new_n293_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT74), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n292_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n604_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n297_), .A2(new_n272_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n601_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n605_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G113gat), .B(G141gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n600_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n608_), .A2(KEYINPUT75), .A3(new_n611_), .A4(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n612_), .A2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n321_), .A2(new_n599_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n554_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n264_), .B1(KEYINPUT99), .B2(KEYINPUT38), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(KEYINPUT99), .A2(KEYINPUT38), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n262_), .A2(new_n621_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n288_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT100), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n316_), .A2(new_n308_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n599_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT101), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n264_), .B1(new_n637_), .B2(new_n554_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n629_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n590_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n623_), .A2(new_n265_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n637_), .A2(new_n642_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G8gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT39), .B(new_n265_), .C1(new_n637_), .C2(new_n642_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1325gat));
  INV_X1    g449(.A(G15gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n402_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n623_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n637_), .A2(new_n652_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n654_), .B2(G15gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n591_), .A2(new_n594_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT104), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n637_), .B2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT42), .Z(new_n664_));
  NAND3_X1  g463(.A1(new_n623_), .A2(new_n659_), .A3(new_n662_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1327gat));
  INV_X1    g465(.A(new_n262_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n289_), .A2(new_n633_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR4_X1   g468(.A1(new_n599_), .A2(new_n667_), .A3(new_n622_), .A4(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n554_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n630_), .A2(new_n289_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n599_), .B2(new_n319_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n595_), .A2(new_n597_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n580_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n491_), .B1(new_n526_), .B2(new_n536_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT98), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT27), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n558_), .B2(new_n492_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n589_), .A3(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n674_), .A2(new_n624_), .A3(new_n675_), .A4(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n561_), .A2(new_n578_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n402_), .A3(new_n660_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT43), .B(new_n319_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n673_), .B1(new_n684_), .B2(KEYINPUT105), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n683_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(new_n319_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n672_), .C1(new_n685_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n684_), .A2(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n689_), .A2(new_n690_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n673_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n697_), .A2(KEYINPUT106), .A3(KEYINPUT44), .A4(new_n672_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n672_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n694_), .A2(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n554_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n671_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n670_), .A2(new_n704_), .A3(new_n642_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n701_), .A2(new_n642_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n704_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT46), .B(new_n706_), .C1(new_n707_), .C2(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  AOI21_X1  g511(.A(G43gat), .B1(new_n670_), .B2(new_n652_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n596_), .A2(G43gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n701_), .B2(new_n714_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n670_), .A2(new_n717_), .A3(new_n662_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n694_), .A2(new_n698_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n660_), .B1(new_n700_), .B2(new_n699_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n721_), .B2(G50gat), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  AOI211_X1 g522(.A(new_n723_), .B(new_n717_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT108), .B(new_n718_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1331gat));
  NOR2_X1   g528(.A1(new_n621_), .A2(new_n288_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n636_), .A2(new_n667_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n554_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n599_), .A2(new_n621_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n262_), .A2(new_n688_), .A3(new_n288_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n735_), .A2(KEYINPUT109), .ZN(new_n736_));
  AOI211_X1 g535(.A(G57gat), .B(new_n624_), .C1(new_n735_), .C2(KEYINPUT109), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n732_), .A2(G57gat), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n731_), .B2(new_n642_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  INV_X1    g541(.A(new_n735_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n740_), .A3(new_n642_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1333gat));
  AOI21_X1  g544(.A(new_n382_), .B1(new_n731_), .B2(new_n652_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n382_), .A3(new_n652_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n731_), .B2(new_n662_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n743_), .A2(new_n751_), .A3(new_n662_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n262_), .A2(new_n669_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n733_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n227_), .A3(new_n554_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n262_), .A2(new_n289_), .A3(new_n621_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n697_), .A2(new_n760_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(new_n554_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n227_), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n228_), .A3(new_n642_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n761_), .A2(new_n642_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n228_), .ZN(G1337gat));
  NAND3_X1  g565(.A1(new_n758_), .A2(new_n222_), .A3(new_n596_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n761_), .A2(new_n652_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n384_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g569(.A1(new_n757_), .A2(G106gat), .A3(new_n660_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n761_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G106gat), .B1(new_n772_), .B2(new_n660_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(KEYINPUT52), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(KEYINPUT52), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n771_), .B(new_n777_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1339gat));
  INV_X1    g580(.A(G113gat), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n622_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n239_), .A2(new_n245_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT12), .B1(new_n212_), .B2(new_n232_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n203_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n246_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT114), .B1(new_n246_), .B2(new_n787_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n246_), .A2(KEYINPUT114), .A3(new_n787_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n788_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n252_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n246_), .A2(KEYINPUT114), .A3(new_n787_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n789_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n794_), .B(new_n251_), .C1(new_n796_), .C2(new_n788_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n793_), .A2(new_n253_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT115), .B1(new_n800_), .B2(new_n616_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n601_), .A2(new_n605_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n609_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(KEYINPUT115), .A3(new_n616_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n803_), .A2(new_n804_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n798_), .A2(new_n799_), .A3(KEYINPUT58), .A4(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n793_), .A2(new_n253_), .A3(new_n797_), .A4(new_n805_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT117), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n808_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT116), .B1(new_n811_), .B2(new_n688_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n319_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n810_), .A2(new_n812_), .A3(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n793_), .A2(new_n621_), .A3(new_n797_), .A4(new_n253_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n805_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT57), .B1(new_n818_), .B2(new_n633_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n634_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n288_), .B1(new_n815_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n621_), .B2(new_n288_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n730_), .A2(KEYINPUT113), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n262_), .A2(new_n319_), .A3(new_n825_), .A4(new_n826_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT54), .Z(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n624_), .B1(new_n823_), .B2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n642_), .A2(new_n597_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT59), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n819_), .A2(new_n821_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n811_), .A2(KEYINPUT116), .A3(new_n688_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n835_), .B2(new_n812_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n828_), .B1(new_n836_), .B2(new_n288_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  INV_X1    g637(.A(new_n831_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n624_), .A4(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n783_), .B1(new_n832_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n811_), .A2(new_n688_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n813_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(new_n834_), .A3(new_n806_), .A4(new_n809_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n289_), .B1(new_n845_), .B2(new_n833_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n554_), .B(new_n831_), .C1(new_n846_), .C2(new_n828_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n842_), .B(new_n782_), .C1(new_n847_), .C2(new_n622_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n823_), .A2(new_n829_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(new_n554_), .A3(new_n621_), .A4(new_n831_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n842_), .B1(new_n851_), .B2(new_n782_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n841_), .B1(new_n849_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT119), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n841_), .B(new_n855_), .C1(new_n849_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1340gat));
  NOR2_X1   g656(.A1(new_n832_), .A2(new_n840_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G120gat), .B1(new_n858_), .B2(new_n262_), .ZN(new_n859_));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n262_), .B2(KEYINPUT60), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(KEYINPUT60), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(KEYINPUT120), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(KEYINPUT120), .B2(new_n861_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n859_), .B1(new_n847_), .B2(new_n864_), .ZN(G1341gat));
  INV_X1    g664(.A(new_n847_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G127gat), .B1(new_n866_), .B2(new_n289_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n858_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n288_), .A2(KEYINPUT121), .ZN(new_n869_));
  MUX2_X1   g668(.A(KEYINPUT121), .B(new_n869_), .S(G127gat), .Z(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n868_), .B2(new_n870_), .ZN(G1342gat));
  OAI21_X1  g670(.A(G134gat), .B1(new_n858_), .B2(new_n319_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n633_), .A2(G134gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n847_), .B2(new_n873_), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n642_), .A2(new_n595_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n830_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n622_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n448_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n262_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n449_), .ZN(G1345gat));
  OR3_X1    g679(.A1(new_n876_), .A2(KEYINPUT122), .A3(new_n288_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n876_), .B2(new_n288_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n876_), .B2(new_n319_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n634_), .A2(new_n444_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n876_), .B2(new_n888_), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n590_), .A2(new_n554_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n652_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n850_), .A2(new_n661_), .A3(new_n893_), .ZN(new_n894_));
  OAI221_X1 g693(.A(G169gat), .B1(KEYINPUT123), .B2(new_n890_), .C1(new_n894_), .C2(new_n622_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n896_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n837_), .A2(new_n662_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n515_), .A2(new_n517_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n621_), .A4(new_n893_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n898_), .A3(new_n901_), .ZN(G1348gat));
  INV_X1    g701(.A(G176gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n894_), .B2(new_n262_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT124), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n850_), .A2(new_n660_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n906_), .A2(new_n903_), .A3(new_n262_), .A4(new_n892_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1349gat));
  NAND4_X1  g707(.A1(new_n850_), .A2(new_n660_), .A3(new_n289_), .A4(new_n893_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n892_), .A2(new_n510_), .A3(new_n288_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n909_), .A2(new_n354_), .B1(new_n899_), .B2(new_n910_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n894_), .B2(new_n319_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n634_), .A2(new_n356_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n894_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1351gat));
  NOR4_X1   g716(.A1(new_n837_), .A2(new_n554_), .A3(new_n590_), .A4(new_n595_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n621_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g719(.A1(new_n918_), .A2(new_n667_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(G204gat), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n428_), .B2(new_n921_), .ZN(G1353gat));
  NAND2_X1  g722(.A1(new_n918_), .A2(new_n289_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n924_), .B2(new_n925_), .ZN(G1354gat));
  NAND2_X1  g727(.A1(new_n918_), .A2(new_n634_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT127), .B(G218gat), .Z(new_n930_));
  NOR2_X1   g729(.A1(new_n319_), .A2(new_n930_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n930_), .B1(new_n918_), .B2(new_n931_), .ZN(G1355gat));
endmodule


