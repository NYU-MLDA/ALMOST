// Benchmark "../Benchmarks/c2670" written by ABC on Fri Feb  4 08:45:06 2022

module c2670  ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241,
    G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253,
    G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269,
    G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452, G483,
    G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384,
    G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066,
    G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106,
    G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193,
    G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205,
    G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240,
    G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252,
    G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268,
    G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452,
    G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348,
    G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996,
    G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105,
    G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474,
    G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_G546_, new_G560_, new_G1385_, new_G157_, new_G547_, new_G258_,
    new_G480_, new_G486_, new_G654_, new_G655_, new_G658_, new_G772_,
    new_G795_, new_G865_, new_G875_, new_G882_, new_G1251_, new_G1254_,
    new_G1261_, new_G1284_, new_G1344_, new_G1351_, new_G1394_, new_G1418_,
    new_G2433_, new_G2434_, new_G2441_, new_G2442_, new_G2449_, new_G2450_,
    new_G2478_, new_G1631_, new_G1655_, new_G1710_, new_G1721_, new_G2682_,
    new_G1955_, new_G1959_, new_G1964_, new_G1969_, new_G1974_, new_G1979_,
    new_G1984_, new_G1989_, new_G1994_, new_G1999_, new_G2001_, new_G2012_,
    new_G2070_, new_G2076_, new_G2082_, new_G2088_, new_G2094_, new_G2099_,
    new_G2103_, new_G2457_, new_G2458_, new_G2461_, new_G2464_, new_G2471_,
    new_G2479_, new_G2482_, new_G2487_, new_G2490_, new_G2495_, new_G2498_,
    new_G2505_, new_G2508_, new_G2675_, new_G2683_, new_G2686_, new_G2691_,
    new_G2694_, new_G2699_, new_G2702_, new_G487_, new_G1475_, new_G1476_,
    new_G1484_, new_G1485_, new_G1493_, new_G1494_, new_G2459_, new_G2460_,
    new_G216_, new_G1253_, new_G1256_, new_G558_, new_G748_, new_G784_,
    new_G807_, new_G821_, new_G825_, new_G829_, new_G833_, new_G837_,
    new_G881_, new_G994_, new_G1273_, new_G1296_, new_G1310_, new_G1314_,
    new_G1318_, new_G1322_, new_G1326_, new_G1406_, new_G1430_, new_G1444_,
    new_G1448_, new_G1452_, new_G1456_, new_G1460_, new_G1477_, new_G1486_,
    new_G1495_, new_G2477_, new_G1499_, new_G2485_, new_G2486_, new_G2493_,
    new_G2494_, new_G1643_, new_G1667_, new_G1681_, new_G1685_, new_G1689_,
    new_G1693_, new_G1697_, new_G1716_, new_G1728_, new_G2681_, new_G1776_,
    new_G2689_, new_G2690_, new_G2697_, new_G2698_, new_G1831_, new_G1893_,
    new_G2007_, new_G2018_, new_G2467_, new_G2468_, new_G2501_, new_G2502_,
    new_G2511_, new_G2512_, new_G2518_, new_G2551_, new_G2559_, new_G2567_,
    new_G2575_, new_G2583_, new_G2591_, new_G2599_, new_G2607_, new_G2615_,
    new_G2623_, new_G2705_, new_G2706_, new_G2735_, new_G2743_, new_G2751_,
    new_G2759_, new_G2767_, new_G2775_, new_G550_, new_G552_, new_G894_,
    new_G1498_, new_G1507_, new_G1508_, new_G1516_, new_G1517_, new_G1775_,
    new_G1784_, new_G1785_, new_G1793_, new_G1794_, new_G2469_, new_G2470_,
    new_G2503_, new_G2504_, new_G2513_, new_G2514_, new_G2707_, new_G2708_,
    new_G551_, new_G553_, new_G818_, new_G819_, new_G820_, new_G822_,
    new_G823_, new_G824_, new_G826_, new_G827_, new_G828_, new_G830_,
    new_G831_, new_G832_, new_G834_, new_G835_, new_G836_, new_G1307_,
    new_G1308_, new_G1309_, new_G1311_, new_G1312_, new_G1313_, new_G1315_,
    new_G1316_, new_G1317_, new_G1319_, new_G1320_, new_G1321_, new_G1323_,
    new_G1324_, new_G1325_, new_G1441_, new_G1442_, new_G1443_, new_G1445_,
    new_G1446_, new_G1447_, new_G1449_, new_G1450_, new_G1451_, new_G1453_,
    new_G1454_, new_G1455_, new_G1457_, new_G1458_, new_G1459_, new_G1481_,
    new_G1490_, new_G1500_, new_G1509_, new_G1518_, new_G1521_, new_G1525_,
    new_G2557_, new_G2565_, new_G2573_, new_G2581_, new_G2589_, new_G2597_,
    new_G2605_, new_G2613_, new_G2621_, new_G2629_, new_G1678_, new_G1679_,
    new_G1680_, new_G1682_, new_G1683_, new_G1684_, new_G1686_, new_G1687_,
    new_G1688_, new_G1690_, new_G1691_, new_G1692_, new_G1694_, new_G1695_,
    new_G1696_, new_G1734_, new_G1736_, new_G1738_, new_G1740_, new_G1742_,
    new_G1744_, new_G1746_, new_G1748_, new_G1750_, new_G1777_, new_G1786_,
    new_G1795_, new_G2023_, new_G2025_, new_G2027_, new_G2029_, new_G2031_,
    new_G2033_, new_G2035_, new_G2037_, new_G2741_, new_G2749_, new_G2757_,
    new_G2765_, new_G2773_, new_G2781_, new_G2515_, new_G2522_, new_G2525_,
    new_G2528_, new_G2730_, new_G554_, new_G838_, new_G841_, new_G846_,
    new_G854_, new_G857_, new_G1327_, new_G1329_, new_G1331_, new_G1333_,
    new_G1335_, new_G1461_, new_G1464_, new_G1467_, new_G1470_, new_G1473_,
    new_G1698_, new_G1701_, new_G1704_, new_G1707_, new_G2634_, new_G1504_,
    new_G1513_, new_G1524_, new_G1528_, new_G1529_, new_G1533_, new_G1538_,
    new_G1541_, new_G1781_, new_G1790_, new_G1806_, new_G1810_, new_G2734_,
    new_G2521_, new_G2524_, new_G2531_, new_G2532_, new_G144_, new_G147_,
    new_G152_, new_G175_, new_G187_, new_G516_, new_G852_, new_G885_,
    new_G887_, new_G893_, new_G1028_, new_G1031_, new_G1035_, new_G1041_,
    new_G1049_, new_G1057_, new_G1060_, new_G1066_, new_G1072_, new_G1078_,
    new_G1213_, new_G1218_, new_G1250_, new_G1387_, new_G1389_, new_G1537_,
    new_G1540_, new_G1735_, new_G1737_, new_G1739_, new_G1741_, new_G1743_,
    new_G1745_, new_G1747_, new_G1749_, new_G1751_, new_G2638_, new_G2024_,
    new_G2026_, new_G2028_, new_G2030_, new_G2032_, new_G2034_, new_G2036_,
    new_G2038_, new_G2154_, new_G2523_, new_G2533_, new_G2534_, new_G2631_,
    new_G2639_, new_G2642_, new_G2647_, new_G2650_, new_G2655_, new_G2658_,
    new_G2665_, new_G2668_, new_G1532_, new_G1536_, new_G1539_, new_G1542_,
    new_G1544_, new_G1547_, new_G2065_, new_G1809_, new_G1813_, new_G1821_,
    new_G1824_, new_G2538_, new_G2546_, new_G2554_, new_G2562_, new_G2570_,
    new_G2578_, new_G2586_, new_G2594_, new_G2602_, new_G2610_, new_G2618_,
    new_G2626_, new_G2738_, new_G2746_, new_G2754_, new_G2762_, new_G2770_,
    new_G2778_, new_G456_, new_G466_, new_G562_, new_G883_, new_G889_,
    new_G891_, new_G1043_, new_G1051_, new_G1062_, new_G1068_, new_G1074_,
    new_G1080_, new_G1225_, new_G1227_, new_G1232_, new_G1234_, new_G1543_,
    new_G1546_, new_G2637_, new_G1753_, new_G2645_, new_G2646_, new_G2653_,
    new_G2654_, new_G1820_, new_G1823_, new_G2107_, new_G2110_, new_G2118_,
    new_G2123_, new_G2151_, new_G2158_, new_G2161_, new_G2164_, new_G2172_,
    new_G2235_, new_G2262_, new_G2350_, new_G2535_, new_G2661_, new_G2662_,
    new_G2671_, new_G2672_, new_G468_, new_G897_, new_G898_, new_G1228_,
    new_G1235_, new_G1545_, new_G1548_, new_G2542_, new_G2550_, new_G1561_,
    new_G2558_, new_G1565_, new_G2566_, new_G1569_, new_G2574_, new_G1573_,
    new_G2582_, new_G1577_, new_G2590_, new_G1581_, new_G2598_, new_G1585_,
    new_G2606_, new_G1589_, new_G2614_, new_G1593_, new_G2622_, new_G1597_,
    new_G2630_, new_G1752_, new_G1761_, new_G1762_, new_G1770_, new_G1771_,
    new_G1822_, new_G1825_, new_G2039_, new_G2742_, new_G2043_, new_G2750_,
    new_G2047_, new_G2758_, new_G2051_, new_G2766_, new_G2055_, new_G2774_,
    new_G2059_, new_G2782_, new_G2663_, new_G2664_, new_G2673_, new_G2674_,
    new_G146_, new_G462_, new_G2113_, new_G2114_, new_G2122_, new_G2129_,
    new_G592_, new_G2167_, new_G2168_, new_G2176_, new_G2241_, new_G2266_,
    new_G743_, new_G749_, new_G886_, new_G995_, new_G1006_, new_G1550_,
    new_G2354_, new_G2541_, new_G1562_, new_G1566_, new_G1570_, new_G1574_,
    new_G1578_, new_G1582_, new_G1586_, new_G1590_, new_G1594_, new_G1598_,
    new_G1754_, new_G1763_, new_G1772_, new_G2040_, new_G2044_, new_G2048_,
    new_G2052_, new_G2056_, new_G2060_, new_G2115_, new_G2126_, new_G2131_,
    new_G2134_, new_G2141_, new_G2144_, new_G2157_, new_G2160_, new_G2169_,
    new_G2177_, new_G2180_, new_G2187_, new_G2190_, new_G2207_, new_G2254_,
    new_G2334_, new_G2342_, new_G2422_, new_G2543_, new_G2709_, new_G2712_,
    new_G2727_, new_G569_, new_G570_, new_G599_, new_G600_, new_G896_,
    new_G1549_, new_G1243_, new_G1245_, new_G1257_, new_G1258_, new_G1563_,
    new_G1567_, new_G1571_, new_G1575_, new_G1579_, new_G1583_, new_G1587_,
    new_G1591_, new_G1595_, new_G1599_, new_G2041_, new_G2045_, new_G2049_,
    new_G2053_, new_G2057_, new_G2061_, new_G2159_, new_G475_, new_G490_,
    new_G496_, new_G502_, new_G508_, new_G765_, new_G769_, new_G571_,
    new_G2121_, new_G579_, new_G587_, new_G2130_, new_G596_, new_G601_,
    new_G2175_, new_G609_, new_G2258_, new_G1014_, new_G1018_, new_G717_,
    new_G723_, new_G729_, new_G735_, new_G753_, new_G2338_, new_G999_,
    new_G1091_, new_G2346_, new_G2426_, new_G1337_, new_G2549_, new_G1552_,
    new_G1600_, new_G1596_, new_G1592_, new_G1588_, new_G1584_, new_G1580_,
    new_G1576_, new_G1572_, new_G1568_, new_G1564_, new_G2062_, new_G2058_,
    new_G2054_, new_G2050_, new_G2046_, new_G2042_, new_G1758_, new_G1767_,
    new_G1798_, new_G1802_, new_G2733_, new_G1829_, new_G2137_, new_G2138_,
    new_G2147_, new_G2148_, new_G2183_, new_G2184_, new_G2193_, new_G2194_,
    new_G2210_, new_G2213_, new_G2715_, new_G2716_, new_G1094_, new_G1096_,
    new_G578_, new_G588_, new_G608_, new_G742_, new_G1005_, new_G1092_,
    new_G1551_, new_G1554_, new_G1555_, new_G1557_, new_G1558_, new_G1828_,
    new_G1845_, new_G1907_, new_G2139_, new_G2140_, new_G2149_, new_G2150_,
    new_G2185_, new_G2186_, new_G2195_, new_G2196_, new_G2717_, new_G2718_,
    new_G154_, new_G155_, new_G763_, new_G767_, new_G531_, new_G537_,
    new_G575_, new_G580_, new_G589_, new_G605_, new_G610_, new_G1012_,
    new_G1016_, new_G705_, new_G711_, new_G1093_, new_G1355_, new_G1553_,
    new_G1556_, new_G1559_, new_G1601_, new_G1801_, new_G1805_, new_G1815_,
    new_G1818_, new_G1830_, new_G1836_, new_G1850_, new_G1898_, new_G1912_,
    new_G2197_, new_G2200_, new_G2214_, new_G2215_, new_G2217_, new_G2220_,
    new_G2722_, new_G492_, new_G498_, new_G504_, new_G510_, new_G519_,
    new_G525_, new_G533_, new_G539_, new_G693_, new_G699_, new_G707_,
    new_G713_, new_G719_, new_G725_, new_G731_, new_G737_, new_G1560_,
    new_G1814_, new_G1817_, new_G2216_, new_G493_, new_G499_, new_G505_,
    new_G511_, new_G521_, new_G527_, new_G534_, new_G540_, new_G584_,
    new_G613_, new_G617_, new_G621_, new_G625_, new_G676_, new_G695_,
    new_G701_, new_G708_, new_G714_, new_G720_, new_G726_, new_G732_,
    new_G738_, new_G1087_, new_G1108_, new_G1361_, new_G1369_, new_G1373_,
    new_G1377_, new_G1607_, new_G1615_, new_G1619_, new_G1623_, new_G1816_,
    new_G1819_, new_G2726_, new_G1842_, new_G1858_, new_G1863_, new_G1866_,
    new_G1868_, new_G1870_, new_G1872_, new_G1874_, new_G1876_, new_G1904_,
    new_G1920_, new_G1925_, new_G1928_, new_G1930_, new_G1932_, new_G1934_,
    new_G1936_, new_G1938_, new_G2203_, new_G2204_, new_G2223_, new_G2224_,
    new_G2238_, new_G522_, new_G528_, new_G696_, new_G702_, new_G1881_,
    new_G1883_, new_G1885_, new_G1887_, new_G1889_, new_G1891_, new_G1943_,
    new_G1945_, new_G1947_, new_G1949_, new_G1951_, new_G1953_, new_G2205_,
    new_G2206_, new_G2225_, new_G2226_, new_G2719_, new_G616_, new_G620_,
    new_G624_, new_G628_, new_G630_, new_G633_, new_G636_, new_G639_,
    new_G645_, new_G2242_, new_G675_, new_G1107_, new_G1368_, new_G1371_,
    new_G1375_, new_G1614_, new_G1617_, new_G1621_, new_G1856_, new_G1861_,
    new_G1918_, new_G1923_, new_G2230_, new_G2246_, new_G2270_, new_G2278_,
    new_G2286_, new_G2294_, new_G2302_, new_G2310_, new_G2358_, new_G2366_,
    new_G2374_, new_G2382_, new_G2390_, new_G2398_, new_G629_, new_G632_,
    new_G635_, new_G638_, new_G646_, new_G677_, new_G1827_, new_G907_,
    new_G915_, new_G922_, new_G924_, new_G937_, new_G946_, new_G1109_,
    new_G1125_, new_G1133_, new_G1140_, new_G1142_, new_G1155_, new_G1164_,
    new_G1378_, new_G1380_, new_G1382_, new_G1624_, new_G1626_, new_G1628_,
    new_G2725_, new_G1859_, new_G1864_, new_G1921_, new_G1926_, new_G2267_,
    new_G2275_, new_G2283_, new_G2291_, new_G2299_, new_G2307_, new_G2318_,
    new_G2326_, new_G2355_, new_G2363_, new_G2371_, new_G2379_, new_G2387_,
    new_G2395_, new_G2406_, new_G2414_, new_G647_, new_G631_, new_G634_,
    new_G637_, new_G640_, new_G2234_, new_G2250_, new_G679_, new_G1826_,
    new_G2274_, new_G2282_, new_G2290_, new_G2298_, new_G2306_, new_G2314_,
    new_G1110_, new_G2362_, new_G2370_, new_G2378_, new_G2386_, new_G2394_,
    new_G2402_, new_G1877_, new_G1879_, new_G1939_, new_G1941_, new_G143_,
    new_G671_, new_G674_, new_G686_, new_G2273_, new_G900_, new_G2281_,
    new_G909_, new_G2289_, new_G917_, new_G2297_, new_G926_, new_G2305_,
    new_G929_, new_G2313_, new_G939_, new_G2322_, new_G2330_, new_G967_,
    new_G1104_, new_G1106_, new_G2361_, new_G1118_, new_G2369_, new_G1127_,
    new_G2377_, new_G1135_, new_G2385_, new_G1144_, new_G2393_, new_G1147_,
    new_G2401_, new_G1157_, new_G2410_, new_G2418_, new_G1184_, new_G2227_,
    new_G2243_, new_G2251_, new_G2259_, new_G2331_, new_G2339_, new_G2347_,
    new_G2419_, new_G687_, new_G899_, new_G908_, new_G916_, new_G925_,
    new_G928_, new_G938_, new_G954_, new_G961_, new_G1117_, new_G1126_,
    new_G1134_, new_G1143_, new_G1146_, new_G1156_, new_G1172_, new_G1179_,
    new_G2315_, new_G2323_, new_G2403_, new_G2411_, new_G2233_, new_G642_,
    new_G2249_, new_G649_, new_G2257_, new_G665_, new_G684_, new_G2265_,
    new_G688_, new_G901_, new_G910_, new_G918_, new_G927_, new_G930_,
    new_G940_, new_G2337_, new_G963_, new_G2345_, new_G1099_, new_G1115_,
    new_G2353_, new_G1119_, new_G1128_, new_G1136_, new_G1145_, new_G1148_,
    new_G1158_, new_G2425_, new_G1181_, new_G641_, new_G648_, new_G664_,
    new_G683_, new_G2321_, new_G948_, new_G2329_, new_G956_, new_G962_,
    new_G1098_, new_G1114_, new_G2409_, new_G1166_, new_G2417_, new_G1174_,
    new_G1180_, new_G643_, new_G650_, new_G666_, new_G681_, new_G690_,
    new_G947_, new_G955_, new_G964_, new_G968_, new_G970_, new_G971_,
    new_G972_, new_G978_, new_G979_, new_G1100_, new_G1112_, new_G1165_,
    new_G1173_, new_G1182_, new_G1185_, new_G1187_, new_G1188_, new_G1189_,
    new_G1195_, new_G1196_, new_G644_, new_G884_, new_G949_, new_G957_,
    new_G969_, new_G973_, new_G1167_, new_G1175_, new_G1186_, new_G1190_,
    new_G680_, new_G682_, new_G895_, new_G1025_, new_G1111_, new_G1113_,
    new_G685_, new_G976_, new_G977_, new_G980_, new_G981_, new_G1116_,
    new_G1193_, new_G1194_, new_G1197_, new_G1198_, new_G982_, new_G983_,
    new_G988_, new_G1027_, new_G1199_, new_G1200_, new_G1205_, new_G984_,
    new_G1085_, new_G1201_, new_G987_, new_G990_, new_G1204_, new_G1207_,
    new_G989_, new_G1206_, new_G991_, new_G1208_, new_G1221_, new_G1238_,
    new_G1239_, new_G1240_, new_G1247_, new_G471_, new_G473_, new_G1088_,
    new_G1089_;
  assign G350 = G452;
  assign G335 = G452;
  assign G409 = G452;
  assign new_G546_ = G1 & G3;
  assign new_G560_ = ~G559;
  assign G369 = G1083;
  assign G367 = G1083;
  assign new_G1385_ = ~G1384;
  assign G411 = G2066;
  assign G337 = G2066;
  assign G384 = G2066;
  assign new_G157_ = G2072 & G2078 & G2090 & G2084;
  assign new_G547_ = ~new_G546_;
  assign G218 = ~G44;
  assign G219 = ~G132;
  assign G220 = ~G82;
  assign G221 = ~G96;
  assign G235 = ~G69;
  assign G236 = ~G120;
  assign G237 = ~G57;
  assign G238 = ~G108;
  assign new_G258_ = G661 & G2 & G15;
  assign new_G480_ = G661;
  assign new_G486_ = G37 & G37;
  assign new_G654_ = G452;
  assign new_G655_ = G8;
  assign new_G658_ = G8;
  assign new_G772_ = G543;
  assign new_G795_ = G651;
  assign new_G865_ = ~G860;
  assign new_G875_ = ~G868;
  assign new_G882_ = G11 & G868;
  assign new_G1251_ = G44 & G96 & G132 & G82;
  assign new_G1254_ = G69 & G108 & G120 & G57;
  assign new_G1261_ = G543;
  assign new_G1284_ = G651;
  assign new_G1344_ = ~G1341;
  assign new_G1351_ = ~G1348;
  assign new_G1394_ = G2104;
  assign new_G1418_ = G2105;
  assign new_G2433_ = ~G2427;
  assign new_G2434_ = ~G2430;
  assign new_G2441_ = ~G2435;
  assign new_G2442_ = ~G2438;
  assign new_G2449_ = ~G2443;
  assign new_G2450_ = ~G2446;
  assign new_G2478_ = ~G2474;
  assign new_G1631_ = G2104;
  assign new_G1655_ = G2105;
  assign new_G1710_ = G16;
  assign new_G1721_ = G16;
  assign new_G2682_ = ~G2678;
  assign new_G1955_ = G7 & G661;
  assign new_G1959_ = ~G1956;
  assign new_G1964_ = ~G1961;
  assign new_G1969_ = ~G1966;
  assign new_G1974_ = ~G1971;
  assign new_G1979_ = ~G1976;
  assign new_G1984_ = ~G1981;
  assign new_G1989_ = ~G1986;
  assign new_G1994_ = ~G1991;
  assign new_G1999_ = ~G1996;
  assign new_G2001_ = G29;
  assign new_G2012_ = G29;
  assign new_G2070_ = ~G2067;
  assign new_G2076_ = ~G2072;
  assign new_G2082_ = ~G2078;
  assign new_G2088_ = ~G2084;
  assign new_G2094_ = ~G2090;
  assign new_G2099_ = ~G2096;
  assign new_G2103_ = ~G2100;
  assign new_G2457_ = ~G2451;
  assign new_G2458_ = ~G2454;
  assign new_G2461_ = G1348;
  assign new_G2464_ = G1341;
  assign new_G2471_ = G1956;
  assign new_G2479_ = G1966;
  assign new_G2482_ = G1961;
  assign new_G2487_ = G1976;
  assign new_G2490_ = G1971;
  assign new_G2495_ = G1986;
  assign new_G2498_ = G1981;
  assign new_G2505_ = G1996;
  assign new_G2508_ = G1991;
  assign new_G2675_ = G2067;
  assign new_G2683_ = G2078;
  assign new_G2686_ = G2072;
  assign new_G2691_ = G2090;
  assign new_G2694_ = G2084;
  assign new_G2699_ = G2100;
  assign new_G2702_ = G2096;
  assign G158 = ~new_G157_;
  assign G259 = ~new_G258_;
  assign new_G487_ = ~new_G486_;
  assign G391 = new_G654_;
  assign new_G1475_ = ~G2430 | ~new_G2433_;
  assign new_G1476_ = ~G2427 | ~new_G2434_;
  assign new_G1484_ = ~G2438 | ~new_G2441_;
  assign new_G1485_ = ~G2435 | ~new_G2442_;
  assign new_G1493_ = ~G2446 | ~new_G2449_;
  assign new_G1494_ = ~G2443 | ~new_G2450_;
  assign new_G2459_ = ~G2454 | ~new_G2457_;
  assign new_G2460_ = ~G2451 | ~new_G2458_;
  assign G173 = G94 & new_G654_;
  assign new_G216_ = G2106 & new_G1955_;
  assign G223 = ~new_G1955_;
  assign G234 = ~G567 | ~new_G1955_;
  assign new_G1253_ = ~new_G1251_;
  assign new_G1256_ = ~new_G1254_;
  assign new_G558_ = new_G1254_ & new_G1251_;
  assign new_G748_ = new_G655_;
  assign new_G784_ = ~new_G772_;
  assign new_G807_ = ~new_G795_;
  assign new_G821_ = new_G795_ & G80 & new_G772_;
  assign new_G825_ = new_G795_ & G68 & new_G772_;
  assign new_G829_ = new_G795_ & G79 & new_G772_;
  assign new_G833_ = new_G795_ & G78 & new_G772_;
  assign new_G837_ = new_G795_ & G77 & new_G772_;
  assign new_G881_ = G11 & new_G875_;
  assign new_G994_ = new_G655_;
  assign new_G1273_ = ~new_G1261_;
  assign new_G1296_ = ~new_G1284_;
  assign new_G1310_ = new_G1284_ & G76 & new_G1261_;
  assign new_G1314_ = new_G1284_ & G75 & new_G1261_;
  assign new_G1318_ = new_G1284_ & G74 & new_G1261_;
  assign new_G1322_ = new_G1284_ & G73 & new_G1261_;
  assign new_G1326_ = new_G1284_ & G72 & new_G1261_;
  assign new_G1406_ = ~new_G1394_;
  assign new_G1430_ = ~new_G1418_;
  assign new_G1444_ = new_G1418_ & G114 & new_G1394_;
  assign new_G1448_ = new_G1418_ & G113 & new_G1394_;
  assign new_G1452_ = new_G1418_ & G112 & new_G1394_;
  assign new_G1456_ = new_G1418_ & G111 & new_G1394_;
  assign new_G1460_ = new_G1394_ & new_G1418_;
  assign new_G1477_ = ~new_G1475_ | ~new_G1476_;
  assign new_G1486_ = ~new_G1484_ | ~new_G1485_;
  assign new_G1495_ = ~new_G1493_ | ~new_G1494_;
  assign new_G2477_ = ~new_G2471_;
  assign new_G1499_ = ~new_G2471_ | ~new_G2478_;
  assign new_G2485_ = ~new_G2479_;
  assign new_G2486_ = ~new_G2482_;
  assign new_G2493_ = ~new_G2487_;
  assign new_G2494_ = ~new_G2490_;
  assign new_G1643_ = ~new_G1631_;
  assign new_G1667_ = ~new_G1655_;
  assign new_G1681_ = new_G1655_ & G118 & new_G1631_;
  assign new_G1685_ = new_G1655_ & G107 & new_G1631_;
  assign new_G1689_ = new_G1655_ & G117 & new_G1631_;
  assign new_G1693_ = new_G1655_ & G116 & new_G1631_;
  assign new_G1697_ = new_G1655_ & G115 & new_G1631_;
  assign new_G1716_ = ~new_G1710_;
  assign new_G1728_ = ~new_G1721_;
  assign new_G2681_ = ~new_G2675_;
  assign new_G1776_ = ~new_G2675_ | ~new_G2682_;
  assign new_G2689_ = ~new_G2683_;
  assign new_G2690_ = ~new_G2686_;
  assign new_G2697_ = ~new_G2691_;
  assign new_G2698_ = ~new_G2694_;
  assign new_G1831_ = new_G658_;
  assign new_G1893_ = new_G658_;
  assign new_G2007_ = ~new_G2001_;
  assign new_G2018_ = ~new_G2012_;
  assign new_G2467_ = ~new_G2461_;
  assign new_G2468_ = ~new_G2464_;
  assign new_G2501_ = ~new_G2495_;
  assign new_G2502_ = ~new_G2498_;
  assign new_G2511_ = ~new_G2505_;
  assign new_G2512_ = ~new_G2508_;
  assign new_G2518_ = ~new_G2459_ | ~new_G2460_;
  assign new_G2551_ = new_G1344_;
  assign new_G2559_ = new_G1351_;
  assign new_G2567_ = new_G1959_;
  assign new_G2575_ = new_G1964_;
  assign new_G2583_ = new_G1969_;
  assign new_G2591_ = new_G1974_;
  assign new_G2599_ = new_G1979_;
  assign new_G2607_ = new_G1984_;
  assign new_G2615_ = new_G1989_;
  assign new_G2623_ = new_G1994_;
  assign new_G2705_ = ~new_G2699_;
  assign new_G2706_ = ~new_G2702_;
  assign new_G2735_ = new_G1999_;
  assign new_G2743_ = new_G2070_;
  assign new_G2751_ = new_G2076_;
  assign new_G2759_ = new_G2082_;
  assign new_G2767_ = new_G2088_;
  assign new_G2775_ = new_G2094_;
  assign G217 = ~new_G216_;
  assign new_G550_ = G2106 & new_G1253_;
  assign new_G552_ = G567 & new_G1256_;
  assign G325 = new_G558_;
  assign new_G894_ = new_G881_ | new_G882_;
  assign new_G1498_ = ~G2474 | ~new_G2477_;
  assign new_G1507_ = ~new_G2482_ | ~new_G2485_;
  assign new_G1508_ = ~new_G2479_ | ~new_G2486_;
  assign new_G1516_ = ~new_G2490_ | ~new_G2493_;
  assign new_G1517_ = ~new_G2487_ | ~new_G2494_;
  assign new_G1775_ = ~G2678 | ~new_G2681_;
  assign new_G1784_ = ~new_G2686_ | ~new_G2689_;
  assign new_G1785_ = ~new_G2683_ | ~new_G2690_;
  assign new_G1793_ = ~new_G2694_ | ~new_G2697_;
  assign new_G1794_ = ~new_G2691_ | ~new_G2698_;
  assign new_G2469_ = ~new_G2464_ | ~new_G2467_;
  assign new_G2470_ = ~new_G2461_ | ~new_G2468_;
  assign new_G2503_ = ~new_G2498_ | ~new_G2501_;
  assign new_G2504_ = ~new_G2495_ | ~new_G2502_;
  assign new_G2513_ = ~new_G2508_ | ~new_G2511_;
  assign new_G2514_ = ~new_G2505_ | ~new_G2512_;
  assign new_G2707_ = ~new_G2702_ | ~new_G2705_;
  assign new_G2708_ = ~new_G2699_ | ~new_G2706_;
  assign G261 = ~new_G558_;
  assign new_G551_ = ~new_G550_;
  assign new_G553_ = ~new_G552_;
  assign new_G818_ = new_G807_ & G93 & new_G784_;
  assign new_G819_ = new_G807_ & G55 & new_G772_;
  assign new_G820_ = new_G795_ & G67 & new_G784_;
  assign new_G822_ = new_G807_ & G81 & new_G784_;
  assign new_G823_ = new_G807_ & G43 & new_G772_;
  assign new_G824_ = new_G795_ & G56 & new_G784_;
  assign new_G826_ = new_G807_ & G92 & new_G784_;
  assign new_G827_ = new_G807_ & G54 & new_G772_;
  assign new_G828_ = new_G795_ & G66 & new_G784_;
  assign new_G830_ = new_G807_ & G91 & new_G784_;
  assign new_G831_ = new_G807_ & G53 & new_G772_;
  assign new_G832_ = new_G795_ & G65 & new_G784_;
  assign new_G834_ = new_G807_ & G90 & new_G784_;
  assign new_G835_ = new_G807_ & G52 & new_G772_;
  assign new_G836_ = new_G795_ & G64 & new_G784_;
  assign new_G1307_ = new_G1296_ & G89 & new_G1273_;
  assign new_G1308_ = new_G1296_ & G51 & new_G1261_;
  assign new_G1309_ = new_G1284_ & G63 & new_G1273_;
  assign new_G1311_ = new_G1296_ & G88 & new_G1273_;
  assign new_G1312_ = new_G1296_ & G50 & new_G1261_;
  assign new_G1313_ = new_G1284_ & G62 & new_G1273_;
  assign new_G1315_ = new_G1296_ & G87 & new_G1273_;
  assign new_G1316_ = new_G1296_ & G49 & new_G1261_;
  assign new_G1317_ = new_G1273_ & new_G1284_;
  assign new_G1319_ = new_G1296_ & G86 & new_G1273_;
  assign new_G1320_ = new_G1296_ & G48 & new_G1261_;
  assign new_G1321_ = new_G1284_ & G61 & new_G1273_;
  assign new_G1323_ = new_G1296_ & G85 & new_G1273_;
  assign new_G1324_ = new_G1296_ & G47 & new_G1261_;
  assign new_G1325_ = new_G1284_ & G60 & new_G1273_;
  assign new_G1441_ = new_G1430_ & G138 & new_G1406_;
  assign new_G1442_ = new_G1430_ & G102 & new_G1394_;
  assign new_G1443_ = new_G1418_ & G126 & new_G1406_;
  assign new_G1445_ = new_G1430_ & G137 & new_G1406_;
  assign new_G1446_ = new_G1430_ & G101 & new_G1394_;
  assign new_G1447_ = new_G1418_ & G125 & new_G1406_;
  assign new_G1449_ = new_G1430_ & G136 & new_G1406_;
  assign new_G1450_ = new_G1430_ & G100 & new_G1394_;
  assign new_G1451_ = new_G1418_ & G124 & new_G1406_;
  assign new_G1453_ = new_G1430_ & G135 & new_G1406_;
  assign new_G1454_ = new_G1430_ & G99 & new_G1394_;
  assign new_G1455_ = new_G1418_ & G123 & new_G1406_;
  assign new_G1457_ = new_G1406_ & new_G1430_;
  assign new_G1458_ = new_G1394_ & new_G1430_;
  assign new_G1459_ = new_G1406_ & new_G1418_;
  assign new_G1481_ = ~new_G1477_;
  assign new_G1490_ = ~new_G1486_;
  assign new_G1500_ = ~new_G1498_ | ~new_G1499_;
  assign new_G1509_ = ~new_G1507_ | ~new_G1508_;
  assign new_G1518_ = ~new_G1516_ | ~new_G1517_;
  assign new_G1521_ = new_G1495_;
  assign new_G1525_ = new_G1495_;
  assign new_G2557_ = ~new_G2551_;
  assign new_G2565_ = ~new_G2559_;
  assign new_G2573_ = ~new_G2567_;
  assign new_G2581_ = ~new_G2575_;
  assign new_G2589_ = ~new_G2583_;
  assign new_G2597_ = ~new_G2591_;
  assign new_G2605_ = ~new_G2599_;
  assign new_G2613_ = ~new_G2607_;
  assign new_G2621_ = ~new_G2615_;
  assign new_G2629_ = ~new_G2623_;
  assign new_G1678_ = new_G1667_ & G142 & new_G1643_;
  assign new_G1679_ = new_G1667_ & G106 & new_G1631_;
  assign new_G1680_ = new_G1655_ & G130 & new_G1643_;
  assign new_G1682_ = new_G1667_ & G131 & new_G1643_;
  assign new_G1683_ = new_G1667_ & G95 & new_G1631_;
  assign new_G1684_ = new_G1655_ & G119 & new_G1643_;
  assign new_G1686_ = new_G1667_ & G141 & new_G1643_;
  assign new_G1687_ = new_G1667_ & G105 & new_G1631_;
  assign new_G1688_ = new_G1655_ & G129 & new_G1643_;
  assign new_G1690_ = new_G1667_ & G140 & new_G1643_;
  assign new_G1691_ = new_G1667_ & G104 & new_G1631_;
  assign new_G1692_ = new_G1655_ & G128 & new_G1643_;
  assign new_G1694_ = new_G1667_ & G139 & new_G1643_;
  assign new_G1695_ = new_G1667_ & G103 & new_G1631_;
  assign new_G1696_ = new_G1655_ & G127 & new_G1643_;
  assign new_G1734_ = G19 & new_G1716_;
  assign new_G1736_ = G4 & new_G1716_;
  assign new_G1738_ = G20 & new_G1716_;
  assign new_G1740_ = G5 & new_G1716_;
  assign new_G1742_ = G21 & new_G1728_;
  assign new_G1744_ = G22 & new_G1728_;
  assign new_G1746_ = G23 & new_G1728_;
  assign new_G1748_ = G6 & new_G1728_;
  assign new_G1750_ = G24 & new_G1728_;
  assign new_G1777_ = ~new_G1775_ | ~new_G1776_;
  assign new_G1786_ = ~new_G1784_ | ~new_G1785_;
  assign new_G1795_ = ~new_G1793_ | ~new_G1794_;
  assign new_G2023_ = G25 & new_G2007_;
  assign new_G2025_ = G32 & new_G2007_;
  assign new_G2027_ = G26 & new_G2007_;
  assign new_G2029_ = G33 & new_G2007_;
  assign new_G2031_ = G27 & new_G2018_;
  assign new_G2033_ = G34 & new_G2018_;
  assign new_G2035_ = G35 & new_G2018_;
  assign new_G2037_ = G28 & new_G2018_;
  assign new_G2741_ = ~new_G2735_;
  assign new_G2749_ = ~new_G2743_;
  assign new_G2757_ = ~new_G2751_;
  assign new_G2765_ = ~new_G2759_;
  assign new_G2773_ = ~new_G2767_;
  assign new_G2781_ = ~new_G2775_;
  assign new_G2515_ = ~new_G2469_ | ~new_G2470_;
  assign new_G2522_ = ~new_G2518_;
  assign new_G2525_ = ~new_G2513_ | ~new_G2514_;
  assign new_G2528_ = ~new_G2503_ | ~new_G2504_;
  assign new_G2730_ = ~new_G2707_ | ~new_G2708_;
  assign new_G554_ = new_G551_ & new_G553_;
  assign new_G838_ = new_G821_ | new_G820_ | new_G818_ | new_G819_;
  assign new_G841_ = new_G825_ | new_G824_ | new_G822_ | new_G823_;
  assign new_G846_ = new_G829_ | new_G828_ | new_G826_ | new_G827_;
  assign new_G854_ = new_G833_ | new_G832_ | new_G830_ | new_G831_;
  assign new_G857_ = new_G837_ | new_G836_ | new_G834_ | new_G835_;
  assign new_G1327_ = new_G1310_ | new_G1309_ | new_G1307_ | new_G1308_;
  assign new_G1329_ = new_G1314_ | new_G1313_ | new_G1311_ | new_G1312_;
  assign new_G1331_ = new_G1318_ | new_G1317_ | new_G1315_ | new_G1316_;
  assign new_G1333_ = new_G1322_ | new_G1321_ | new_G1319_ | new_G1320_;
  assign new_G1335_ = new_G1326_ | new_G1325_ | new_G1323_ | new_G1324_;
  assign new_G1461_ = new_G1444_ | new_G1443_ | new_G1441_ | new_G1442_;
  assign new_G1464_ = new_G1448_ | new_G1447_ | new_G1445_ | new_G1446_;
  assign new_G1467_ = new_G1452_ | new_G1451_ | new_G1449_ | new_G1450_;
  assign new_G1470_ = new_G1456_ | new_G1455_ | new_G1453_ | new_G1454_;
  assign new_G1473_ = new_G1460_ | new_G1459_ | new_G1457_ | new_G1458_;
  assign new_G1698_ = new_G1685_ | new_G1684_ | new_G1682_ | new_G1683_;
  assign new_G1701_ = new_G1689_ | new_G1688_ | new_G1686_ | new_G1687_;
  assign new_G1704_ = new_G1693_ | new_G1692_ | new_G1690_ | new_G1691_;
  assign new_G1707_ = new_G1697_ | new_G1696_ | new_G1694_ | new_G1695_;
  assign new_G2634_ = new_G1681_ | new_G1680_ | new_G1678_ | new_G1679_;
  assign G319 = new_G554_;
  assign new_G1504_ = ~new_G1500_;
  assign new_G1513_ = ~new_G1509_;
  assign new_G1524_ = ~new_G1521_;
  assign new_G1528_ = ~new_G1525_;
  assign new_G1529_ = new_G1518_;
  assign new_G1533_ = new_G1518_;
  assign new_G1538_ = new_G1521_ & new_G1486_ & new_G1477_;
  assign new_G1541_ = new_G1525_ & new_G1490_ & new_G1481_;
  assign new_G1781_ = ~new_G1777_;
  assign new_G1790_ = ~new_G1786_;
  assign new_G1806_ = new_G1795_;
  assign new_G1810_ = new_G1795_;
  assign new_G2734_ = ~new_G2730_;
  assign new_G2521_ = ~new_G2515_;
  assign new_G2524_ = ~new_G2515_ | ~new_G2522_;
  assign new_G2531_ = ~new_G2525_;
  assign new_G2532_ = ~new_G2528_;
  assign new_G144_ = new_G838_ & G860;
  assign new_G147_ = new_G846_ & G860;
  assign new_G152_ = new_G841_ & G860;
  assign G160 = ~new_G1464_;
  assign G162 = ~new_G1467_;
  assign G164 = ~new_G1461_;
  assign G166 = ~new_G1329_;
  assign G168 = ~new_G1327_;
  assign G171 = ~new_G857_;
  assign new_G175_ = new_G554_ & G36 & new_G480_ & G483;
  assign new_G187_ = new_G547_ & new_G554_ & new_G480_ & G483;
  assign new_G516_ = new_G838_;
  assign new_G852_ = ~new_G846_;
  assign new_G885_ = new_G841_ & new_G875_;
  assign new_G887_ = new_G846_ & new_G875_;
  assign new_G893_ = new_G1327_ & G868;
  assign new_G1028_ = ~new_G838_;
  assign new_G1031_ = ~new_G841_;
  assign new_G1035_ = ~new_G846_;
  assign new_G1041_ = new_G854_;
  assign new_G1049_ = new_G857_;
  assign new_G1057_ = new_G1327_;
  assign new_G1060_ = new_G1329_;
  assign new_G1066_ = new_G1331_;
  assign new_G1072_ = new_G1333_;
  assign new_G1078_ = new_G1335_;
  assign new_G1213_ = ~new_G2099_ | ~new_G1470_;
  assign new_G1218_ = ~new_G2103_ | ~new_G1473_;
  assign new_G1250_ = new_G1704_;
  assign new_G1387_ = new_G1461_ & new_G1385_;
  assign new_G1389_ = ~new_G1464_;
  assign new_G1537_ = new_G1524_ & new_G1481_ & new_G1486_;
  assign new_G1540_ = new_G1528_ & new_G1477_ & new_G1490_;
  assign new_G1735_ = new_G841_ & new_G1710_;
  assign new_G1737_ = new_G846_ & new_G1710_;
  assign new_G1739_ = new_G854_ & new_G1710_;
  assign new_G1741_ = new_G857_ & new_G1710_;
  assign new_G1743_ = new_G1327_ & new_G1721_;
  assign new_G1745_ = new_G1329_ & new_G1721_;
  assign new_G1747_ = new_G1331_ & new_G1721_;
  assign new_G1749_ = new_G1333_ & new_G1721_;
  assign new_G1751_ = new_G1335_ & new_G1721_;
  assign new_G2638_ = ~new_G2634_;
  assign new_G2024_ = new_G1698_ & new_G2001_;
  assign new_G2026_ = new_G1701_ & new_G2001_;
  assign new_G2028_ = new_G1704_ & new_G2001_;
  assign new_G2030_ = new_G1707_ & new_G2001_;
  assign new_G2032_ = new_G1461_ & new_G2012_;
  assign new_G2034_ = new_G1464_ & new_G2012_;
  assign new_G2036_ = new_G1467_ & new_G2012_;
  assign new_G2038_ = new_G1470_ & new_G2012_;
  assign new_G2154_ = new_G841_;
  assign new_G2523_ = ~new_G2518_ | ~new_G2521_;
  assign new_G2533_ = ~new_G2528_ | ~new_G2531_;
  assign new_G2534_ = ~new_G2525_ | ~new_G2532_;
  assign new_G2631_ = new_G1698_;
  assign new_G2639_ = new_G1704_;
  assign new_G2642_ = new_G1701_;
  assign new_G2647_ = new_G1461_;
  assign new_G2650_ = new_G1707_;
  assign new_G2655_ = new_G1467_;
  assign new_G2658_ = new_G1464_;
  assign new_G2665_ = new_G1473_;
  assign new_G2668_ = new_G1470_;
  assign G153 = new_G865_ | new_G152_;
  assign G176 = ~new_G175_;
  assign G188 = ~new_G187_;
  assign G299 = new_G1041_;
  assign G301 = new_G1049_;
  assign G286 = new_G1057_;
  assign G303 = new_G1060_;
  assign G288 = new_G1066_;
  assign G305 = new_G1072_;
  assign G290 = new_G1078_;
  assign new_G1532_ = ~new_G1529_;
  assign new_G1536_ = ~new_G1533_;
  assign new_G1539_ = ~new_G1537_ & ~new_G1538_;
  assign new_G1542_ = ~new_G1540_ & ~new_G1541_;
  assign new_G1544_ = new_G1529_ & new_G1509_ & new_G1500_;
  assign new_G1547_ = new_G1533_ & new_G1513_ & new_G1504_;
  assign new_G2065_ = new_G2037_ | new_G2038_;
  assign new_G1809_ = ~new_G1806_;
  assign new_G1813_ = ~new_G1810_;
  assign new_G1821_ = new_G1806_ & new_G1786_ & new_G1777_;
  assign new_G1824_ = new_G1810_ & new_G1790_ & new_G1781_;
  assign new_G2538_ = ~new_G2523_ | ~new_G2524_;
  assign new_G2546_ = ~new_G2533_ | ~new_G2534_;
  assign new_G2554_ = new_G1734_ | new_G1735_;
  assign new_G2562_ = new_G1736_ | new_G1737_;
  assign new_G2570_ = new_G1738_ | new_G1739_;
  assign new_G2578_ = new_G1740_ | new_G1741_;
  assign new_G2586_ = new_G1742_ | new_G1743_;
  assign new_G2594_ = new_G1744_ | new_G1745_;
  assign new_G2602_ = new_G1746_ | new_G1747_;
  assign new_G2610_ = new_G1748_ | new_G1749_;
  assign new_G2618_ = new_G1750_ | new_G1751_;
  assign new_G2626_ = new_G2023_ | new_G2024_;
  assign new_G2738_ = new_G2025_ | new_G2026_;
  assign new_G2746_ = new_G2027_ | new_G2028_;
  assign new_G2754_ = new_G2029_ | new_G2030_;
  assign new_G2762_ = new_G2031_ | new_G2032_;
  assign new_G2770_ = new_G2033_ | new_G2034_;
  assign new_G2778_ = new_G2035_ | new_G2036_;
  assign new_G456_ = G40 & new_G1389_ & new_G1387_;
  assign new_G466_ = ~new_G1387_;
  assign new_G562_ = ~new_G560_ | ~new_G852_;
  assign new_G883_ = new_G516_ & new_G875_;
  assign new_G889_ = new_G1049_ & G868;
  assign new_G891_ = new_G1041_ & new_G875_;
  assign new_G1043_ = ~new_G1041_;
  assign new_G1051_ = ~new_G1049_;
  assign new_G1062_ = ~new_G1060_;
  assign new_G1068_ = ~new_G1066_;
  assign new_G1074_ = ~new_G1072_;
  assign new_G1080_ = ~new_G1078_;
  assign new_G1225_ = new_G2099_ & new_G1213_;
  assign new_G1227_ = new_G1213_ & new_G1470_;
  assign new_G1232_ = new_G2103_ & new_G1218_;
  assign new_G1234_ = new_G1218_ & new_G1473_;
  assign new_G1543_ = new_G1532_ & new_G1504_ & new_G1509_;
  assign new_G1546_ = new_G1536_ & new_G1500_ & new_G1513_;
  assign new_G2637_ = ~new_G2631_;
  assign new_G1753_ = ~new_G2631_ | ~new_G2638_;
  assign new_G2645_ = ~new_G2639_;
  assign new_G2646_ = ~new_G2642_;
  assign new_G2653_ = ~new_G2647_;
  assign new_G2654_ = ~new_G2650_;
  assign new_G1820_ = new_G1809_ & new_G1781_ & new_G1786_;
  assign new_G1823_ = new_G1813_ & new_G1777_ & new_G1790_;
  assign new_G2107_ = new_G1031_;
  assign new_G2110_ = new_G1028_;
  assign new_G2118_ = new_G1035_;
  assign new_G2123_ = ~new_G1057_;
  assign new_G2151_ = ~new_G852_;
  assign new_G2158_ = ~new_G2154_;
  assign new_G2161_ = new_G1031_;
  assign new_G2164_ = new_G1028_;
  assign new_G2172_ = new_G1035_;
  assign new_G2235_ = new_G516_;
  assign new_G2262_ = new_G1035_;
  assign new_G2350_ = new_G1035_;
  assign new_G2535_ = ~new_G1542_ | ~new_G1539_;
  assign new_G2661_ = ~new_G2655_;
  assign new_G2662_ = ~new_G2658_;
  assign new_G2671_ = ~new_G2665_;
  assign new_G2672_ = ~new_G2668_;
  assign new_G468_ = new_G466_ & G40 & new_G1389_;
  assign new_G897_ = new_G887_ | new_G889_;
  assign new_G898_ = new_G891_ | new_G893_;
  assign new_G1228_ = new_G1225_ | new_G1227_;
  assign new_G1235_ = new_G1232_ | new_G1234_;
  assign new_G1545_ = ~new_G1543_ & ~new_G1544_;
  assign new_G1548_ = ~new_G1546_ & ~new_G1547_;
  assign new_G2542_ = ~new_G2538_;
  assign new_G2550_ = ~new_G2546_;
  assign new_G1561_ = ~new_G2554_ | ~new_G2557_;
  assign new_G2558_ = ~new_G2554_;
  assign new_G1565_ = ~new_G2562_ | ~new_G2565_;
  assign new_G2566_ = ~new_G2562_;
  assign new_G1569_ = ~new_G2570_ | ~new_G2573_;
  assign new_G2574_ = ~new_G2570_;
  assign new_G1573_ = ~new_G2578_ | ~new_G2581_;
  assign new_G2582_ = ~new_G2578_;
  assign new_G1577_ = ~new_G2586_ | ~new_G2589_;
  assign new_G2590_ = ~new_G2586_;
  assign new_G1581_ = ~new_G2594_ | ~new_G2597_;
  assign new_G2598_ = ~new_G2594_;
  assign new_G1585_ = ~new_G2602_ | ~new_G2605_;
  assign new_G2606_ = ~new_G2602_;
  assign new_G1589_ = ~new_G2610_ | ~new_G2613_;
  assign new_G2614_ = ~new_G2610_;
  assign new_G1593_ = ~new_G2618_ | ~new_G2621_;
  assign new_G2622_ = ~new_G2618_;
  assign new_G1597_ = ~new_G2626_ | ~new_G2629_;
  assign new_G2630_ = ~new_G2626_;
  assign new_G1752_ = ~new_G2634_ | ~new_G2637_;
  assign new_G1761_ = ~new_G2642_ | ~new_G2645_;
  assign new_G1762_ = ~new_G2639_ | ~new_G2646_;
  assign new_G1770_ = ~new_G2650_ | ~new_G2653_;
  assign new_G1771_ = ~new_G2647_ | ~new_G2654_;
  assign new_G1822_ = ~new_G1820_ & ~new_G1821_;
  assign new_G1825_ = ~new_G1823_ & ~new_G1824_;
  assign new_G2039_ = ~new_G2738_ | ~new_G2741_;
  assign new_G2742_ = ~new_G2738_;
  assign new_G2043_ = ~new_G2746_ | ~new_G2749_;
  assign new_G2750_ = ~new_G2746_;
  assign new_G2047_ = ~new_G2754_ | ~new_G2757_;
  assign new_G2758_ = ~new_G2754_;
  assign new_G2051_ = ~new_G2762_ | ~new_G2765_;
  assign new_G2766_ = ~new_G2762_;
  assign new_G2055_ = ~new_G2770_ | ~new_G2773_;
  assign new_G2774_ = ~new_G2770_;
  assign new_G2059_ = ~new_G2778_ | ~new_G2781_;
  assign new_G2782_ = ~new_G2778_;
  assign new_G2663_ = ~new_G2658_ | ~new_G2661_;
  assign new_G2664_ = ~new_G2655_ | ~new_G2662_;
  assign new_G2673_ = ~new_G2668_ | ~new_G2671_;
  assign new_G2674_ = ~new_G2665_ | ~new_G2672_;
  assign new_G146_ = new_G562_ & new_G865_;
  assign new_G462_ = ~new_G456_;
  assign new_G2113_ = ~new_G2107_;
  assign new_G2114_ = ~new_G2110_;
  assign new_G2122_ = ~new_G2118_;
  assign new_G2129_ = ~new_G2123_;
  assign new_G592_ = new_G562_;
  assign new_G2167_ = ~new_G2161_;
  assign new_G2168_ = ~new_G2164_;
  assign new_G2176_ = ~new_G2172_;
  assign new_G2241_ = ~new_G2235_;
  assign new_G2266_ = ~new_G2262_;
  assign new_G743_ = ~new_G456_;
  assign new_G749_ = new_G456_;
  assign new_G886_ = new_G562_ & G868;
  assign G284 = new_G897_;
  assign G321 = new_G897_;
  assign G297 = new_G898_;
  assign G280 = new_G898_;
  assign new_G995_ = new_G456_;
  assign new_G1006_ = ~new_G456_;
  assign new_G1550_ = ~new_G2535_ | ~new_G2542_;
  assign new_G2354_ = ~new_G2350_;
  assign new_G2541_ = ~new_G2535_;
  assign new_G1562_ = ~new_G2551_ | ~new_G2558_;
  assign new_G1566_ = ~new_G2559_ | ~new_G2566_;
  assign new_G1570_ = ~new_G2567_ | ~new_G2574_;
  assign new_G1574_ = ~new_G2575_ | ~new_G2582_;
  assign new_G1578_ = ~new_G2583_ | ~new_G2590_;
  assign new_G1582_ = ~new_G2591_ | ~new_G2598_;
  assign new_G1586_ = ~new_G2599_ | ~new_G2606_;
  assign new_G1590_ = ~new_G2607_ | ~new_G2614_;
  assign new_G1594_ = ~new_G2615_ | ~new_G2622_;
  assign new_G1598_ = ~new_G2623_ | ~new_G2630_;
  assign new_G1754_ = ~new_G1752_ | ~new_G1753_;
  assign new_G1763_ = ~new_G1761_ | ~new_G1762_;
  assign new_G1772_ = ~new_G1770_ | ~new_G1771_;
  assign new_G2040_ = ~new_G2735_ | ~new_G2742_;
  assign new_G2044_ = ~new_G2743_ | ~new_G2750_;
  assign new_G2048_ = ~new_G2751_ | ~new_G2758_;
  assign new_G2052_ = ~new_G2759_ | ~new_G2766_;
  assign new_G2056_ = ~new_G2767_ | ~new_G2774_;
  assign new_G2060_ = ~new_G2775_ | ~new_G2782_;
  assign new_G2115_ = new_G1043_;
  assign new_G2126_ = new_G1051_;
  assign new_G2131_ = new_G1068_;
  assign new_G2134_ = new_G1062_;
  assign new_G2141_ = new_G1080_;
  assign new_G2144_ = new_G1074_;
  assign new_G2157_ = ~new_G2151_;
  assign new_G2160_ = ~new_G2151_ | ~new_G2158_;
  assign new_G2169_ = new_G1043_;
  assign new_G2177_ = new_G1068_;
  assign new_G2180_ = new_G1062_;
  assign new_G2187_ = new_G1080_;
  assign new_G2190_ = new_G1074_;
  assign new_G2207_ = ~new_G562_;
  assign new_G2254_ = new_G1043_;
  assign new_G2334_ = new_G1051_;
  assign new_G2342_ = new_G1043_;
  assign new_G2422_ = new_G1051_;
  assign new_G2543_ = ~new_G1548_ | ~new_G1545_;
  assign new_G2709_ = ~new_G2673_ | ~new_G2674_;
  assign new_G2712_ = ~new_G2663_ | ~new_G2664_;
  assign new_G2727_ = ~new_G1825_ | ~new_G1822_;
  assign G148 = new_G146_ | new_G147_;
  assign new_G569_ = ~new_G2110_ | ~new_G2113_;
  assign new_G570_ = ~new_G2107_ | ~new_G2114_;
  assign new_G599_ = ~new_G2164_ | ~new_G2167_;
  assign new_G600_ = ~new_G2161_ | ~new_G2168_;
  assign new_G896_ = new_G885_ | new_G886_;
  assign new_G1549_ = ~new_G2538_ | ~new_G2541_;
  assign new_G1243_ = ~new_G1228_;
  assign new_G1245_ = ~new_G1235_;
  assign new_G1257_ = new_G468_;
  assign new_G1258_ = new_G468_;
  assign new_G1563_ = ~new_G1561_ | ~new_G1562_;
  assign new_G1567_ = ~new_G1565_ | ~new_G1566_;
  assign new_G1571_ = ~new_G1569_ | ~new_G1570_;
  assign new_G1575_ = ~new_G1573_ | ~new_G1574_;
  assign new_G1579_ = ~new_G1577_ | ~new_G1578_;
  assign new_G1583_ = ~new_G1581_ | ~new_G1582_;
  assign new_G1587_ = ~new_G1585_ | ~new_G1586_;
  assign new_G1591_ = ~new_G1589_ | ~new_G1590_;
  assign new_G1595_ = ~new_G1593_ | ~new_G1594_;
  assign new_G1599_ = ~new_G1597_ | ~new_G1598_;
  assign new_G2041_ = ~new_G2039_ | ~new_G2040_;
  assign new_G2045_ = ~new_G2043_ | ~new_G2044_;
  assign new_G2049_ = ~new_G2047_ | ~new_G2048_;
  assign new_G2053_ = ~new_G2051_ | ~new_G2052_;
  assign new_G2057_ = ~new_G2055_ | ~new_G2056_;
  assign new_G2061_ = ~new_G2059_ | ~new_G2060_;
  assign new_G2159_ = ~new_G2154_ | ~new_G2157_;
  assign new_G475_ = new_G462_;
  assign new_G490_ = new_G1078_ & new_G743_;
  assign new_G496_ = new_G1698_ & new_G743_;
  assign new_G502_ = new_G1701_ & new_G743_;
  assign new_G508_ = new_G1250_ & new_G743_;
  assign new_G765_ = new_G1057_ & new_G749_;
  assign new_G769_ = new_G1060_ & new_G749_;
  assign new_G571_ = ~new_G569_ | ~new_G570_;
  assign new_G2121_ = ~new_G2115_;
  assign new_G579_ = ~new_G2115_ | ~new_G2122_;
  assign new_G587_ = ~new_G2126_ | ~new_G2129_;
  assign new_G2130_ = ~new_G2126_;
  assign new_G596_ = ~new_G592_;
  assign new_G601_ = ~new_G599_ | ~new_G600_;
  assign new_G2175_ = ~new_G2169_;
  assign new_G609_ = ~new_G2169_ | ~new_G2176_;
  assign new_G2258_ = ~new_G2254_;
  assign new_G1014_ = new_G1057_ & new_G995_;
  assign new_G1018_ = new_G1060_ & new_G995_;
  assign new_G717_ = new_G1078_ & new_G1006_;
  assign new_G723_ = new_G1698_ & new_G1006_;
  assign new_G729_ = new_G1701_ & new_G1006_;
  assign new_G735_ = new_G1250_ & new_G1006_;
  assign new_G753_ = ~new_G749_;
  assign G282 = new_G896_;
  assign G323 = new_G896_;
  assign new_G2338_ = ~new_G2334_;
  assign new_G999_ = ~new_G995_;
  assign new_G1091_ = ~new_G1549_ | ~new_G1550_;
  assign new_G2346_ = ~new_G2342_;
  assign new_G2426_ = ~new_G2422_;
  assign new_G1337_ = new_G462_;
  assign new_G2549_ = ~new_G2543_;
  assign new_G1552_ = ~new_G2543_ | ~new_G2550_;
  assign new_G1600_ = ~new_G1599_;
  assign new_G1596_ = ~new_G1595_;
  assign new_G1592_ = ~new_G1591_;
  assign new_G1588_ = ~new_G1587_;
  assign new_G1584_ = ~new_G1583_;
  assign new_G1580_ = ~new_G1579_;
  assign new_G1576_ = ~new_G1575_;
  assign new_G1572_ = ~new_G1571_;
  assign new_G1568_ = ~new_G1567_;
  assign new_G1564_ = ~new_G1563_;
  assign new_G2062_ = ~new_G2061_;
  assign new_G2058_ = ~new_G2057_;
  assign new_G2054_ = ~new_G2053_;
  assign new_G2050_ = ~new_G2049_;
  assign new_G2046_ = ~new_G2045_;
  assign new_G2042_ = ~new_G2041_;
  assign new_G1758_ = ~new_G1754_;
  assign new_G1767_ = ~new_G1763_;
  assign new_G1798_ = new_G1772_;
  assign new_G1802_ = new_G1772_;
  assign new_G2733_ = ~new_G2727_;
  assign new_G1829_ = ~new_G2727_ | ~new_G2734_;
  assign new_G2137_ = ~new_G2131_;
  assign new_G2138_ = ~new_G2134_;
  assign new_G2147_ = ~new_G2141_;
  assign new_G2148_ = ~new_G2144_;
  assign new_G2183_ = ~new_G2177_;
  assign new_G2184_ = ~new_G2180_;
  assign new_G2193_ = ~new_G2187_;
  assign new_G2194_ = ~new_G2190_;
  assign new_G2210_ = ~new_G2159_ | ~new_G2160_;
  assign new_G2213_ = ~new_G2207_;
  assign new_G2715_ = ~new_G2709_;
  assign new_G2716_ = ~new_G2712_;
  assign new_G1094_ = new_G1235_ & new_G1245_;
  assign new_G1096_ = new_G1228_ & new_G1243_;
  assign new_G578_ = ~new_G2118_ | ~new_G2121_;
  assign new_G588_ = ~new_G2123_ | ~new_G2130_;
  assign new_G608_ = ~new_G2172_ | ~new_G2175_;
  assign new_G742_ = new_G1257_;
  assign new_G1005_ = new_G1257_;
  assign new_G1092_ = ~new_G1091_;
  assign new_G1551_ = ~new_G2546_ | ~new_G2549_;
  assign new_G1554_ = new_G1584_ & new_G1588_ & new_G1592_ & new_G1600_ & new_G1596_;
  assign new_G1555_ = new_G1564_ & new_G1568_ & new_G1572_ & new_G1580_ & new_G1576_;
  assign new_G1557_ = new_G2065_ & new_G2062_;
  assign new_G1558_ = new_G2042_ & new_G2046_ & new_G2050_ & new_G2058_ & new_G2054_;
  assign new_G1828_ = ~new_G2730_ | ~new_G2733_;
  assign new_G1845_ = new_G1258_;
  assign new_G1907_ = new_G1258_;
  assign new_G2139_ = ~new_G2134_ | ~new_G2137_;
  assign new_G2140_ = ~new_G2131_ | ~new_G2138_;
  assign new_G2149_ = ~new_G2144_ | ~new_G2147_;
  assign new_G2150_ = ~new_G2141_ | ~new_G2148_;
  assign new_G2185_ = ~new_G2180_ | ~new_G2183_;
  assign new_G2186_ = ~new_G2177_ | ~new_G2184_;
  assign new_G2195_ = ~new_G2190_ | ~new_G2193_;
  assign new_G2196_ = ~new_G2187_ | ~new_G2194_;
  assign new_G2717_ = ~new_G2712_ | ~new_G2715_;
  assign new_G2718_ = ~new_G2709_ | ~new_G2716_;
  assign new_G154_ = new_G1094_ | new_G1245_;
  assign new_G155_ = new_G1096_ | new_G1243_;
  assign new_G763_ = new_G1057_ & new_G753_;
  assign new_G767_ = new_G1060_ & new_G753_;
  assign new_G531_ = new_G1066_ & new_G753_;
  assign new_G537_ = new_G1072_ & new_G753_;
  assign new_G575_ = ~new_G571_;
  assign new_G580_ = ~new_G578_ | ~new_G579_;
  assign new_G589_ = ~new_G587_ | ~new_G588_;
  assign new_G605_ = ~new_G601_;
  assign new_G610_ = ~new_G608_ | ~new_G609_;
  assign new_G1012_ = new_G1057_ & new_G999_;
  assign new_G1016_ = new_G1060_ & new_G999_;
  assign new_G705_ = new_G1066_ & new_G999_;
  assign new_G711_ = new_G1072_ & new_G999_;
  assign new_G1093_ = new_G1092_ & G14;
  assign new_G1355_ = new_G475_;
  assign new_G1553_ = ~new_G1551_ | ~new_G1552_;
  assign new_G1556_ = new_G1554_ & new_G1555_;
  assign new_G1559_ = new_G1557_ & new_G1558_;
  assign new_G1601_ = new_G1337_;
  assign new_G1801_ = ~new_G1798_;
  assign new_G1805_ = ~new_G1802_;
  assign new_G1815_ = new_G1798_ & new_G1763_ & new_G1754_;
  assign new_G1818_ = new_G1802_ & new_G1767_ & new_G1758_;
  assign new_G1830_ = ~new_G1828_ | ~new_G1829_;
  assign new_G1836_ = new_G475_;
  assign new_G1850_ = new_G475_;
  assign new_G1898_ = new_G1337_;
  assign new_G1912_ = new_G1337_;
  assign new_G2197_ = ~new_G2149_ | ~new_G2150_;
  assign new_G2200_ = ~new_G2139_ | ~new_G2140_;
  assign new_G2214_ = ~new_G2210_;
  assign new_G2215_ = ~new_G2210_ | ~new_G2213_;
  assign new_G2217_ = ~new_G2195_ | ~new_G2196_;
  assign new_G2220_ = ~new_G2185_ | ~new_G2186_;
  assign new_G2722_ = ~new_G2717_ | ~new_G2718_;
  assign G156 = ~new_G154_ | ~new_G155_;
  assign new_G492_ = new_G490_ & new_G742_;
  assign new_G498_ = new_G496_ & new_G742_;
  assign new_G504_ = new_G502_ & new_G742_;
  assign new_G510_ = new_G508_ & new_G742_;
  assign new_G519_ = new_G763_ | new_G765_;
  assign new_G525_ = new_G767_ | new_G769_;
  assign new_G533_ = new_G531_ & new_G748_;
  assign new_G539_ = new_G537_ & new_G748_;
  assign new_G693_ = new_G1012_ | new_G1014_;
  assign new_G699_ = new_G1016_ | new_G1018_;
  assign new_G707_ = new_G705_ & new_G994_;
  assign new_G713_ = new_G711_ & new_G994_;
  assign new_G719_ = new_G717_ & new_G1005_;
  assign new_G725_ = new_G723_ & new_G1005_;
  assign new_G731_ = new_G729_ & new_G1005_;
  assign new_G737_ = new_G735_ & new_G1005_;
  assign G401 = new_G1093_;
  assign new_G1560_ = new_G894_ & new_G1556_ & new_G1559_;
  assign new_G1814_ = new_G1801_ & new_G1758_ & new_G1763_;
  assign new_G1817_ = new_G1805_ & new_G1754_ & new_G1767_;
  assign new_G2216_ = ~new_G2207_ | ~new_G2214_;
  assign G227 = ~new_G1830_;
  assign G229 = ~new_G1553_;
  assign new_G493_ = ~new_G492_;
  assign new_G499_ = ~new_G498_;
  assign new_G505_ = ~new_G504_;
  assign new_G511_ = ~new_G510_;
  assign new_G521_ = new_G519_ & new_G748_;
  assign new_G527_ = new_G525_ & new_G748_;
  assign new_G534_ = ~new_G533_;
  assign new_G540_ = ~new_G539_;
  assign new_G584_ = ~new_G580_;
  assign new_G613_ = new_G589_;
  assign new_G617_ = new_G589_;
  assign new_G621_ = new_G610_;
  assign new_G625_ = new_G610_;
  assign new_G676_ = new_G1344_ & new_G1355_;
  assign new_G695_ = new_G693_ & new_G994_;
  assign new_G701_ = new_G699_ & new_G994_;
  assign new_G708_ = ~new_G707_;
  assign new_G714_ = ~new_G713_;
  assign new_G720_ = ~new_G719_;
  assign new_G726_ = ~new_G725_;
  assign new_G732_ = ~new_G731_;
  assign new_G738_ = ~new_G737_;
  assign new_G1087_ = ~new_G1093_;
  assign new_G1108_ = new_G1344_ & new_G1601_;
  assign new_G1361_ = ~new_G1355_;
  assign new_G1369_ = new_G1351_ & new_G1355_;
  assign new_G1373_ = new_G1959_ & new_G1355_;
  assign new_G1377_ = new_G1964_ & new_G1355_;
  assign G311 = new_G1560_;
  assign new_G1607_ = ~new_G1601_;
  assign new_G1615_ = new_G1351_ & new_G1601_;
  assign new_G1619_ = new_G1959_ & new_G1601_;
  assign new_G1623_ = new_G1964_ & new_G1601_;
  assign new_G1816_ = ~new_G1814_ & ~new_G1815_;
  assign new_G1819_ = ~new_G1817_ & ~new_G1818_;
  assign new_G2726_ = ~new_G2722_;
  assign new_G1842_ = ~new_G1836_;
  assign new_G1858_ = new_G1969_ & new_G1836_;
  assign new_G1863_ = new_G1974_ & new_G1836_;
  assign new_G1866_ = new_G1979_ & new_G1836_;
  assign new_G1868_ = new_G1984_ & new_G1836_;
  assign new_G1870_ = new_G1989_ & new_G1850_;
  assign new_G1872_ = new_G1994_ & new_G1850_;
  assign new_G1874_ = new_G1999_ & new_G1850_;
  assign new_G1876_ = new_G2070_ & new_G1850_;
  assign new_G1904_ = ~new_G1898_;
  assign new_G1920_ = new_G1969_ & new_G1898_;
  assign new_G1925_ = new_G1974_ & new_G1898_;
  assign new_G1928_ = new_G1979_ & new_G1898_;
  assign new_G1930_ = new_G1984_ & new_G1898_;
  assign new_G1932_ = new_G1989_ & new_G1912_;
  assign new_G1934_ = new_G1994_ & new_G1912_;
  assign new_G1936_ = new_G1999_ & new_G1912_;
  assign new_G1938_ = new_G2070_ & new_G1912_;
  assign new_G2203_ = ~new_G2197_;
  assign new_G2204_ = ~new_G2200_;
  assign new_G2223_ = ~new_G2217_;
  assign new_G2224_ = ~new_G2220_;
  assign new_G2238_ = ~new_G2215_ | ~new_G2216_;
  assign G150 = ~new_G1560_;
  assign new_G522_ = ~new_G521_;
  assign new_G528_ = ~new_G527_;
  assign new_G696_ = ~new_G695_;
  assign new_G702_ = ~new_G701_;
  assign new_G1881_ = new_G1866_ & new_G1831_;
  assign new_G1883_ = new_G1868_ & new_G1831_;
  assign new_G1885_ = new_G1870_ & new_G1845_;
  assign new_G1887_ = new_G1872_ & new_G1845_;
  assign new_G1889_ = new_G1874_ & new_G1845_;
  assign new_G1891_ = new_G1876_ & new_G1845_;
  assign new_G1943_ = new_G1928_ & new_G1893_;
  assign new_G1945_ = new_G1930_ & new_G1893_;
  assign new_G1947_ = new_G1932_ & new_G1907_;
  assign new_G1949_ = new_G1934_ & new_G1907_;
  assign new_G1951_ = new_G1936_ & new_G1907_;
  assign new_G1953_ = new_G1938_ & new_G1907_;
  assign new_G2205_ = ~new_G2200_ | ~new_G2203_;
  assign new_G2206_ = ~new_G2197_ | ~new_G2204_;
  assign new_G2225_ = ~new_G2220_ | ~new_G2223_;
  assign new_G2226_ = ~new_G2217_ | ~new_G2224_;
  assign new_G2719_ = ~new_G1819_ | ~new_G1816_;
  assign new_G616_ = ~new_G613_;
  assign new_G620_ = ~new_G617_;
  assign new_G624_ = ~new_G621_;
  assign new_G628_ = ~new_G625_;
  assign new_G630_ = new_G613_ & new_G580_ & new_G571_;
  assign new_G633_ = new_G617_ & new_G584_ & new_G575_;
  assign new_G636_ = new_G621_ & new_G601_ & new_G592_;
  assign new_G639_ = new_G625_ & new_G605_ & new_G596_;
  assign new_G645_ = ~new_G2238_ | ~new_G2241_;
  assign new_G2242_ = ~new_G2238_;
  assign new_G675_ = new_G1999_ & new_G1361_;
  assign new_G1107_ = new_G1999_ & new_G1607_;
  assign new_G1368_ = new_G2070_ & new_G1361_;
  assign new_G1371_ = new_G2076_ & new_G1361_;
  assign new_G1375_ = new_G2082_ & new_G1361_;
  assign new_G1614_ = new_G2070_ & new_G1607_;
  assign new_G1617_ = new_G2076_ & new_G1607_;
  assign new_G1621_ = new_G2082_ & new_G1607_;
  assign new_G1856_ = new_G2088_ & new_G1842_;
  assign new_G1861_ = new_G2094_ & new_G1842_;
  assign new_G1918_ = new_G2088_ & new_G1904_;
  assign new_G1923_ = new_G2094_ & new_G1904_;
  assign new_G2230_ = ~new_G2205_ | ~new_G2206_;
  assign new_G2246_ = ~new_G2225_ | ~new_G2226_;
  assign new_G2270_ = new_G511_;
  assign new_G2278_ = new_G505_;
  assign new_G2286_ = new_G499_;
  assign new_G2294_ = new_G493_;
  assign new_G2302_ = new_G540_;
  assign new_G2310_ = new_G534_;
  assign new_G2358_ = new_G738_;
  assign new_G2366_ = new_G732_;
  assign new_G2374_ = new_G726_;
  assign new_G2382_ = new_G720_;
  assign new_G2390_ = new_G714_;
  assign new_G2398_ = new_G708_;
  assign new_G629_ = new_G616_ & new_G575_ & new_G580_;
  assign new_G632_ = new_G620_ & new_G571_ & new_G584_;
  assign new_G635_ = new_G624_ & new_G596_ & new_G601_;
  assign new_G638_ = new_G628_ & new_G592_ & new_G605_;
  assign new_G646_ = ~new_G2235_ | ~new_G2242_;
  assign new_G677_ = new_G675_ | new_G676_;
  assign new_G1827_ = ~new_G2719_ | ~new_G2726_;
  assign new_G907_ = new_G1891_ & new_G511_;
  assign new_G915_ = new_G1889_ & new_G505_;
  assign new_G922_ = new_G1887_ & new_G499_;
  assign new_G924_ = new_G493_ & new_G1885_;
  assign new_G937_ = new_G1883_ & new_G540_;
  assign new_G946_ = new_G1881_ & new_G534_;
  assign new_G1109_ = new_G1107_ | new_G1108_;
  assign new_G1125_ = new_G1953_ & new_G738_;
  assign new_G1133_ = new_G1951_ & new_G732_;
  assign new_G1140_ = new_G1949_ & new_G726_;
  assign new_G1142_ = new_G720_ & new_G1947_;
  assign new_G1155_ = new_G1945_ & new_G714_;
  assign new_G1164_ = new_G1943_ & new_G708_;
  assign new_G1378_ = new_G1368_ | new_G1369_;
  assign new_G1380_ = new_G1371_ | new_G1373_;
  assign new_G1382_ = new_G1375_ | new_G1377_;
  assign new_G1624_ = new_G1614_ | new_G1615_;
  assign new_G1626_ = new_G1617_ | new_G1619_;
  assign new_G1628_ = new_G1621_ | new_G1623_;
  assign new_G2725_ = ~new_G2719_;
  assign new_G1859_ = new_G1856_ | new_G1858_;
  assign new_G1864_ = new_G1861_ | new_G1863_;
  assign new_G1921_ = new_G1918_ | new_G1920_;
  assign new_G1926_ = new_G1923_ | new_G1925_;
  assign new_G2267_ = new_G1891_;
  assign new_G2275_ = new_G1889_;
  assign new_G2283_ = new_G1887_;
  assign new_G2291_ = new_G1885_;
  assign new_G2299_ = new_G1883_;
  assign new_G2307_ = new_G1881_;
  assign new_G2318_ = new_G528_;
  assign new_G2326_ = new_G522_;
  assign new_G2355_ = new_G1953_;
  assign new_G2363_ = new_G1951_;
  assign new_G2371_ = new_G1949_;
  assign new_G2379_ = new_G1947_;
  assign new_G2387_ = new_G1945_;
  assign new_G2395_ = new_G1943_;
  assign new_G2406_ = new_G702_;
  assign new_G2414_ = new_G696_;
  assign new_G647_ = ~new_G645_ | ~new_G646_;
  assign new_G631_ = ~new_G629_ & ~new_G630_;
  assign new_G634_ = ~new_G632_ & ~new_G633_;
  assign new_G637_ = ~new_G635_ & ~new_G636_;
  assign new_G640_ = ~new_G638_ & ~new_G639_;
  assign new_G2234_ = ~new_G2230_;
  assign new_G2250_ = ~new_G2246_;
  assign new_G679_ = new_G677_ & new_G1031_;
  assign new_G1826_ = ~new_G2722_ | ~new_G2725_;
  assign new_G2274_ = ~new_G2270_;
  assign new_G2282_ = ~new_G2278_;
  assign new_G2290_ = ~new_G2286_;
  assign new_G2298_ = ~new_G2294_;
  assign new_G2306_ = ~new_G2302_;
  assign new_G2314_ = ~new_G2310_;
  assign new_G1110_ = new_G1109_ & new_G1031_;
  assign new_G2362_ = ~new_G2358_;
  assign new_G2370_ = ~new_G2366_;
  assign new_G2378_ = ~new_G2374_;
  assign new_G2386_ = ~new_G2382_;
  assign new_G2394_ = ~new_G2390_;
  assign new_G2402_ = ~new_G2398_;
  assign new_G1877_ = new_G1859_ & new_G1831_;
  assign new_G1879_ = new_G1864_ & new_G1831_;
  assign new_G1939_ = new_G1921_ & new_G1893_;
  assign new_G1941_ = new_G1926_ & new_G1893_;
  assign new_G143_ = new_G647_ & new_G865_;
  assign new_G671_ = new_G1380_ & new_G1043_;
  assign new_G674_ = new_G1378_ & new_G1035_;
  assign new_G686_ = ~new_G1826_ | ~new_G1827_;
  assign new_G2273_ = ~new_G2267_;
  assign new_G900_ = ~new_G2267_ | ~new_G2274_;
  assign new_G2281_ = ~new_G2275_;
  assign new_G909_ = ~new_G2275_ | ~new_G2282_;
  assign new_G2289_ = ~new_G2283_;
  assign new_G917_ = ~new_G2283_ | ~new_G2290_;
  assign new_G2297_ = ~new_G2291_;
  assign new_G926_ = ~new_G2291_ | ~new_G2298_;
  assign new_G2305_ = ~new_G2299_;
  assign new_G929_ = ~new_G2299_ | ~new_G2306_;
  assign new_G2313_ = ~new_G2307_;
  assign new_G939_ = ~new_G2307_ | ~new_G2314_;
  assign new_G2322_ = ~new_G2318_;
  assign new_G2330_ = ~new_G2326_;
  assign new_G967_ = new_G1382_ & new_G1051_;
  assign new_G1104_ = new_G1626_ & new_G1043_;
  assign new_G1106_ = new_G1624_ & new_G1035_;
  assign new_G2361_ = ~new_G2355_;
  assign new_G1118_ = ~new_G2355_ | ~new_G2362_;
  assign new_G2369_ = ~new_G2363_;
  assign new_G1127_ = ~new_G2363_ | ~new_G2370_;
  assign new_G2377_ = ~new_G2371_;
  assign new_G1135_ = ~new_G2371_ | ~new_G2378_;
  assign new_G2385_ = ~new_G2379_;
  assign new_G1144_ = ~new_G2379_ | ~new_G2386_;
  assign new_G2393_ = ~new_G2387_;
  assign new_G1147_ = ~new_G2387_ | ~new_G2394_;
  assign new_G2401_ = ~new_G2395_;
  assign new_G1157_ = ~new_G2395_ | ~new_G2402_;
  assign new_G2410_ = ~new_G2406_;
  assign new_G2418_ = ~new_G2414_;
  assign new_G1184_ = new_G1628_ & new_G1051_;
  assign new_G2227_ = ~new_G634_ | ~new_G631_;
  assign new_G2243_ = ~new_G640_ | ~new_G637_;
  assign new_G2251_ = new_G1380_;
  assign new_G2259_ = new_G1378_;
  assign new_G2331_ = new_G1382_;
  assign new_G2339_ = new_G1626_;
  assign new_G2347_ = new_G1624_;
  assign new_G2419_ = new_G1628_;
  assign G145 = new_G143_ | new_G144_;
  assign new_G687_ = ~new_G686_;
  assign new_G899_ = ~new_G2270_ | ~new_G2273_;
  assign new_G908_ = ~new_G2278_ | ~new_G2281_;
  assign new_G916_ = ~new_G2286_ | ~new_G2289_;
  assign new_G925_ = ~new_G2294_ | ~new_G2297_;
  assign new_G928_ = ~new_G2302_ | ~new_G2305_;
  assign new_G938_ = ~new_G2310_ | ~new_G2313_;
  assign new_G954_ = new_G1879_ & new_G528_;
  assign new_G961_ = new_G1877_ & new_G522_;
  assign new_G1117_ = ~new_G2358_ | ~new_G2361_;
  assign new_G1126_ = ~new_G2366_ | ~new_G2369_;
  assign new_G1134_ = ~new_G2374_ | ~new_G2377_;
  assign new_G1143_ = ~new_G2382_ | ~new_G2385_;
  assign new_G1146_ = ~new_G2390_ | ~new_G2393_;
  assign new_G1156_ = ~new_G2398_ | ~new_G2401_;
  assign new_G1172_ = new_G1941_ & new_G702_;
  assign new_G1179_ = new_G1939_ & new_G696_;
  assign new_G2315_ = new_G1879_;
  assign new_G2323_ = new_G1877_;
  assign new_G2403_ = new_G1941_;
  assign new_G2411_ = new_G1939_;
  assign new_G2233_ = ~new_G2227_;
  assign new_G642_ = ~new_G2227_ | ~new_G2234_;
  assign new_G2249_ = ~new_G2243_;
  assign new_G649_ = ~new_G2243_ | ~new_G2250_;
  assign new_G2257_ = ~new_G2251_;
  assign new_G665_ = ~new_G2251_ | ~new_G2258_;
  assign new_G684_ = ~new_G2259_ | ~new_G2266_;
  assign new_G2265_ = ~new_G2259_;
  assign new_G688_ = new_G687_ & new_G487_;
  assign new_G901_ = ~new_G899_ | ~new_G900_;
  assign new_G910_ = ~new_G908_ | ~new_G909_;
  assign new_G918_ = ~new_G916_ | ~new_G917_;
  assign new_G927_ = ~new_G925_ | ~new_G926_;
  assign new_G930_ = ~new_G928_ | ~new_G929_;
  assign new_G940_ = ~new_G938_ | ~new_G939_;
  assign new_G2337_ = ~new_G2331_;
  assign new_G963_ = ~new_G2331_ | ~new_G2338_;
  assign new_G2345_ = ~new_G2339_;
  assign new_G1099_ = ~new_G2339_ | ~new_G2346_;
  assign new_G1115_ = ~new_G2347_ | ~new_G2354_;
  assign new_G2353_ = ~new_G2347_;
  assign new_G1119_ = ~new_G1117_ | ~new_G1118_;
  assign new_G1128_ = ~new_G1126_ | ~new_G1127_;
  assign new_G1136_ = ~new_G1134_ | ~new_G1135_;
  assign new_G1145_ = ~new_G1143_ | ~new_G1144_;
  assign new_G1148_ = ~new_G1146_ | ~new_G1147_;
  assign new_G1158_ = ~new_G1156_ | ~new_G1157_;
  assign new_G2425_ = ~new_G2419_;
  assign new_G1181_ = ~new_G2419_ | ~new_G2426_;
  assign new_G641_ = ~new_G2230_ | ~new_G2233_;
  assign new_G648_ = ~new_G2246_ | ~new_G2249_;
  assign new_G664_ = ~new_G2254_ | ~new_G2257_;
  assign new_G683_ = ~new_G2262_ | ~new_G2265_;
  assign G395 = new_G688_;
  assign new_G2321_ = ~new_G2315_;
  assign new_G948_ = ~new_G2315_ | ~new_G2322_;
  assign new_G2329_ = ~new_G2323_;
  assign new_G956_ = ~new_G2323_ | ~new_G2330_;
  assign new_G962_ = ~new_G2334_ | ~new_G2337_;
  assign new_G1098_ = ~new_G2342_ | ~new_G2345_;
  assign new_G1114_ = ~new_G2350_ | ~new_G2353_;
  assign new_G2409_ = ~new_G2403_;
  assign new_G1166_ = ~new_G2403_ | ~new_G2410_;
  assign new_G2417_ = ~new_G2411_;
  assign new_G1174_ = ~new_G2411_ | ~new_G2418_;
  assign new_G1180_ = ~new_G2422_ | ~new_G2425_;
  assign new_G643_ = ~new_G641_ | ~new_G642_;
  assign new_G650_ = ~new_G648_ | ~new_G649_;
  assign new_G666_ = ~new_G664_ | ~new_G665_;
  assign new_G681_ = ~new_G683_ | ~new_G684_;
  assign new_G690_ = ~new_G688_;
  assign new_G947_ = ~new_G2318_ | ~new_G2321_;
  assign new_G955_ = ~new_G2326_ | ~new_G2329_;
  assign new_G964_ = ~new_G962_ | ~new_G963_;
  assign new_G968_ = new_G901_ & new_G918_ & new_G910_ & new_G927_;
  assign new_G970_ = new_G901_ & new_G915_;
  assign new_G971_ = new_G922_ & new_G910_ & new_G901_;
  assign new_G972_ = new_G910_ & new_G924_ & new_G918_ & new_G901_;
  assign new_G978_ = new_G930_ & new_G946_;
  assign new_G979_ = new_G954_ & new_G940_ & new_G930_;
  assign new_G1100_ = ~new_G1098_ | ~new_G1099_;
  assign new_G1112_ = ~new_G1114_ | ~new_G1115_;
  assign new_G1165_ = ~new_G2406_ | ~new_G2409_;
  assign new_G1173_ = ~new_G2414_ | ~new_G2417_;
  assign new_G1182_ = ~new_G1180_ | ~new_G1181_;
  assign new_G1185_ = new_G1119_ & new_G1136_ & new_G1128_ & new_G1145_;
  assign new_G1187_ = new_G1119_ & new_G1133_;
  assign new_G1188_ = new_G1140_ & new_G1128_ & new_G1119_;
  assign new_G1189_ = new_G1128_ & new_G1142_ & new_G1136_ & new_G1119_;
  assign new_G1195_ = new_G1148_ & new_G1164_;
  assign new_G1196_ = new_G1172_ & new_G1158_ & new_G1148_;
  assign new_G644_ = ~new_G643_;
  assign new_G884_ = new_G650_ & G868;
  assign new_G949_ = ~new_G947_ | ~new_G948_;
  assign new_G957_ = ~new_G955_ | ~new_G956_;
  assign new_G969_ = ~new_G968_;
  assign new_G973_ = new_G972_ | new_G971_ | new_G907_ | new_G970_;
  assign new_G1167_ = ~new_G1165_ | ~new_G1166_;
  assign new_G1175_ = ~new_G1173_ | ~new_G1174_;
  assign new_G1186_ = ~new_G1185_;
  assign new_G1190_ = new_G1189_ | new_G1188_ | new_G1125_ | new_G1187_;
  assign new_G680_ = new_G666_ & new_G674_;
  assign new_G682_ = new_G679_ & new_G681_ & new_G666_;
  assign new_G895_ = new_G883_ | new_G884_;
  assign new_G1025_ = new_G644_ & new_G487_;
  assign new_G1111_ = new_G1100_ & new_G1106_;
  assign new_G1113_ = new_G1110_ & new_G1112_ & new_G1100_;
  assign new_G685_ = new_G682_ | new_G671_ | new_G680_;
  assign G295 = new_G895_;
  assign G331 = new_G895_;
  assign new_G976_ = ~new_G973_;
  assign new_G977_ = new_G957_ & new_G930_ & new_G949_ & new_G940_ & new_G964_;
  assign new_G980_ = new_G940_ & new_G961_ & new_G949_ & new_G930_;
  assign new_G981_ = new_G940_ & new_G967_ & new_G930_ & new_G957_ & new_G949_;
  assign G397 = new_G1025_;
  assign new_G1116_ = new_G1113_ | new_G1104_ | new_G1111_;
  assign new_G1193_ = ~new_G1190_;
  assign new_G1194_ = new_G1175_ & new_G1148_ & new_G1167_ & new_G1158_ & new_G1182_;
  assign new_G1197_ = new_G1158_ & new_G1179_ & new_G1167_ & new_G1148_;
  assign new_G1198_ = new_G1158_ & new_G1184_ & new_G1148_ & new_G1175_ & new_G1167_;
  assign new_G982_ = new_G981_ | new_G980_ | new_G979_ | new_G937_ | new_G978_;
  assign new_G983_ = new_G977_ & new_G685_;
  assign new_G988_ = ~new_G976_ | ~new_G969_;
  assign new_G1027_ = ~new_G1025_;
  assign new_G1199_ = new_G1198_ | new_G1197_ | new_G1196_ | new_G1155_ | new_G1195_;
  assign new_G1200_ = new_G1194_ & new_G1116_;
  assign new_G1205_ = ~new_G1193_ | ~new_G1186_;
  assign new_G984_ = new_G982_ | new_G983_;
  assign new_G1085_ = new_G1830_ & new_G690_ & new_G1027_;
  assign new_G1201_ = new_G1199_ | new_G1200_;
  assign new_G987_ = ~new_G984_;
  assign new_G990_ = new_G988_ & new_G984_;
  assign new_G1204_ = ~new_G1201_;
  assign new_G1207_ = new_G1205_ & new_G1201_;
  assign new_G989_ = new_G973_ & new_G987_;
  assign new_G1206_ = new_G1190_ & new_G1204_;
  assign new_G991_ = new_G989_ | new_G990_;
  assign new_G1208_ = new_G1206_ | new_G1207_;
  assign G329 = new_G1208_;
  assign new_G1221_ = ~new_G1208_ | ~new_G991_;
  assign new_G1238_ = new_G1208_ & new_G1221_;
  assign new_G1239_ = new_G1221_ & new_G991_;
  assign new_G1240_ = new_G1238_ | new_G1239_;
  assign new_G1247_ = ~new_G1240_;
  assign new_G471_ = new_G1240_ & new_G1247_;
  assign new_G473_ = new_G471_ | new_G1247_;
  assign G231 = ~new_G473_;
  assign new_G1088_ = new_G473_ & new_G1553_ & new_G1087_;
  assign new_G1089_ = new_G554_ & new_G1085_ & new_G1088_;
  assign G308 = new_G1089_;
  assign G225 = ~new_G1089_;
endmodule


