//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  XNOR2_X1  g000(.A(KEYINPUT26), .B(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(G183gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n206_));
  OAI21_X1  g005(.A(G183gat), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT81), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT81), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n204_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT83), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT82), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n210_), .A2(new_n211_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n211_), .B1(new_n210_), .B2(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n219_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT23), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n221_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n212_), .B(KEYINPUT83), .Z(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n231_), .B(new_n232_), .C1(G176gat), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT30), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT86), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT30), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT86), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  INV_X1    g043(.A(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT85), .B(G15gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n250_), .B1(new_n237_), .B2(KEYINPUT86), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G127gat), .B(G134gat), .Z(new_n254_));
  XOR2_X1   g053(.A(G113gat), .B(G120gat), .Z(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT31), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(new_n253_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n250_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n261_), .B2(new_n252_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n266_), .B2(KEYINPUT92), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT90), .B(G204gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(G197gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n264_), .B1(G197gat), .B2(G204gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n269_), .B2(G197gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT91), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n265_), .B1(new_n270_), .B2(KEYINPUT21), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G228gat), .A2(G233gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT87), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  INV_X1    g085(.A(G141gat), .ZN(new_n287_));
  INV_X1    g086(.A(G148gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n289_), .B(new_n290_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n282_), .B1(new_n285_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n281_), .B1(new_n280_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n295_), .B2(new_n280_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n287_), .A2(new_n288_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT88), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n278_), .B(new_n279_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n278_), .A2(KEYINPUT93), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT93), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(new_n273_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n307_), .A2(new_n309_), .B1(KEYINPUT29), .B2(new_n300_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n306_), .B1(new_n310_), .B2(new_n279_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT95), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n306_), .B(KEYINPUT95), .C1(new_n310_), .C2(new_n279_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n314_), .B(KEYINPUT94), .Z(new_n317_));
  OAI211_X1 g116(.A(new_n306_), .B(new_n317_), .C1(new_n310_), .C2(new_n279_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT96), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n304_), .A2(new_n305_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G22gat), .B(G50gat), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n304_), .A2(new_n305_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n323_), .A2(new_n327_), .A3(new_n325_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT96), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n318_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n316_), .A2(new_n320_), .A3(new_n331_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n329_), .A2(new_n330_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n317_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n311_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n337_), .B2(new_n319_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n278_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n227_), .B2(new_n235_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT19), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n345_), .A2(new_n202_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT24), .A4(new_n212_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n225_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT97), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n348_), .A2(new_n349_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n232_), .A2(KEYINPUT98), .B1(new_n225_), .B2(new_n230_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT98), .ZN(new_n353_));
  INV_X1    g152(.A(G176gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n213_), .A2(new_n353_), .B1(new_n354_), .B2(new_n233_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n352_), .A2(KEYINPUT99), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT99), .B1(new_n352_), .B2(new_n355_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n350_), .B(new_n351_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT20), .B(new_n344_), .C1(new_n358_), .C2(new_n278_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n341_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n227_), .A2(new_n340_), .A3(new_n235_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT20), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n358_), .B2(new_n278_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n344_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n301_), .A2(new_n303_), .A3(new_n256_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n300_), .A2(new_n256_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n373_), .B(new_n376_), .C1(new_n379_), .C2(new_n375_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G29gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G85gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT0), .B(G57gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n372_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n371_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n352_), .A2(new_n355_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n391_), .A2(new_n348_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n307_), .A2(new_n309_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT100), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n236_), .A2(new_n278_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n393_), .B2(KEYINPUT20), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n343_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT101), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT101), .B(new_n343_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n361_), .A2(new_n363_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(new_n343_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n370_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n390_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n364_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n341_), .A2(new_n359_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n369_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n369_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n384_), .B1(new_n379_), .B2(new_n373_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n375_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n375_), .B2(new_n374_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n416_), .B2(new_n373_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n411_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n380_), .A2(new_n386_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n384_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT33), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n389_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n339_), .B1(new_n408_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(new_n413_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT27), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n387_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT102), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n411_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n365_), .A2(KEYINPUT102), .A3(new_n369_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT27), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n404_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n369_), .B1(new_n436_), .B2(new_n402_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n428_), .B(new_n430_), .C1(new_n435_), .C2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n263_), .B1(new_n425_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n429_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n257_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n261_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n339_), .B(new_n428_), .C1(new_n435_), .C2(new_n437_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT76), .B(G15gat), .ZN(new_n449_));
  INV_X1    g248(.A(G22gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(KEYINPUT76), .A2(G15gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT76), .A2(G15gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(G22gat), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT14), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT77), .B(G1gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(G8gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n448_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n455_), .A2(new_n458_), .A3(new_n448_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G29gat), .B(G36gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT79), .ZN(new_n467_));
  INV_X1    g266(.A(new_n465_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n469_), .B2(KEYINPUT78), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n451_), .A2(new_n454_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n458_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n447_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n465_), .B1(new_n473_), .B2(new_n459_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT79), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n466_), .B1(new_n470_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n469_), .A2(KEYINPUT78), .A3(new_n467_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT79), .B1(new_n474_), .B2(new_n475_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n462_), .A4(new_n465_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n479_), .A3(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n465_), .B(KEYINPUT15), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n462_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n478_), .A3(new_n469_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n446_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT66), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  NAND3_X1  g305(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n499_), .A2(new_n502_), .A3(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT67), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G85gat), .ZN(new_n513_));
  INV_X1    g312(.A(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT8), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT68), .B1(new_n509_), .B2(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n512_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n499_), .A2(new_n502_), .A3(new_n508_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NOR4_X1   g324(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n512_), .A2(new_n518_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT8), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n517_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n531_));
  NOR2_X1   g330(.A1(new_n510_), .A2(new_n511_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT10), .B(G99gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT64), .B(G106gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n502_), .A2(new_n508_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n484_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  OAI221_X1 g343(.A(new_n541_), .B1(KEYINPUT35), .B2(new_n544_), .C1(new_n465_), .C2(new_n540_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT35), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n547_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n551_), .A2(new_n556_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n548_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n559_), .A2(new_n552_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n495_), .B(new_n557_), .C1(new_n558_), .C2(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n552_), .A2(new_n559_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT37), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G120gat), .B(G148gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT72), .ZN(new_n567_));
  XOR2_X1   g366(.A(G176gat), .B(G204gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G71gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT69), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(G71gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(G78gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT69), .B(G71gat), .ZN(new_n580_));
  INV_X1    g379(.A(G78gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT11), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n582_), .A3(KEYINPUT11), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n579_), .A2(new_n582_), .A3(KEYINPUT11), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n529_), .A2(new_n591_), .A3(new_n539_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n591_), .B1(new_n529_), .B2(new_n539_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n573_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT70), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n597_), .B(new_n573_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n588_), .A2(new_n590_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n524_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n499_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n512_), .A2(new_n518_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n519_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n601_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n600_), .B1(new_n606_), .B2(new_n538_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(KEYINPUT12), .A3(new_n592_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n540_), .A2(new_n609_), .A3(new_n600_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n573_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n571_), .B1(new_n599_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n599_), .A2(new_n611_), .A3(new_n571_), .ZN(new_n614_));
  OAI22_X1  g413(.A1(new_n613_), .A2(new_n614_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n612_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G231gat), .ZN(new_n621_));
  INV_X1    g420(.A(G233gat), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n600_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n462_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n623_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n623_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n591_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n462_), .B1(new_n630_), .B2(new_n626_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT17), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT17), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n628_), .A2(new_n631_), .A3(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n565_), .A2(new_n620_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n494_), .A2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(new_n440_), .A3(new_n457_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT38), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT38), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n562_), .A2(new_n563_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n446_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n493_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n619_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n643_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n440_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n647_), .A2(new_n648_), .A3(new_n656_), .ZN(G1324gat));
  NAND2_X1  g456(.A1(new_n406_), .A2(new_n412_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n427_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n658_), .A2(new_n659_), .B1(new_n427_), .B2(new_n426_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G8gat), .B1(new_n655_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT39), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n645_), .A2(G8gat), .A3(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g464(.A(new_n263_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n645_), .A2(G15gat), .A3(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT103), .Z(new_n668_));
  OAI21_X1  g467(.A(G15gat), .B1(new_n655_), .B2(new_n666_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT41), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(KEYINPUT41), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n670_), .A3(new_n671_), .ZN(G1326gat));
  OAI21_X1  g471(.A(G22gat), .B1(new_n655_), .B2(new_n339_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT42), .ZN(new_n674_));
  INV_X1    g473(.A(new_n339_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n450_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT104), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n645_), .B2(new_n677_), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n650_), .A2(new_n643_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n620_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n494_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n494_), .A2(KEYINPUT105), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n429_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n561_), .A2(new_n564_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n446_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(new_n565_), .C1(new_n439_), .C2(new_n445_), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n642_), .B(new_n653_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT44), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(G29gat), .A3(new_n429_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n691_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n695_), .A2(new_n652_), .A3(new_n619_), .A4(new_n643_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n687_), .B1(new_n694_), .B2(new_n698_), .ZN(G1328gat));
  XOR2_X1   g498(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n660_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n698_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n660_), .A2(G36gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n683_), .A2(new_n684_), .A3(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n683_), .A2(new_n684_), .A3(new_n704_), .A4(new_n706_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n700_), .B1(new_n703_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT108), .B(new_n700_), .C1(new_n703_), .C2(new_n710_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n703_), .A2(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT46), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n713_), .A2(new_n714_), .A3(new_n716_), .ZN(G1329gat));
  OAI21_X1  g516(.A(new_n245_), .B1(new_n685_), .B2(new_n666_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n693_), .A2(G43gat), .A3(new_n263_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n698_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n686_), .B2(new_n675_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n693_), .A2(G50gat), .A3(new_n675_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n698_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n446_), .A2(new_n652_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n726_), .A2(new_n620_), .A3(new_n642_), .A4(new_n688_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G57gat), .B1(new_n728_), .B2(new_n429_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n483_), .A2(new_n486_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n489_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n642_), .A3(new_n490_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n619_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n651_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n440_), .A2(KEYINPUT109), .ZN(new_n737_));
  MUX2_X1   g536(.A(KEYINPUT109), .B(new_n737_), .S(G57gat), .Z(new_n738_));
  AOI21_X1  g537(.A(new_n729_), .B1(new_n736_), .B2(new_n738_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n735_), .B2(new_n660_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT48), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n660_), .A2(G64gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n727_), .B2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n735_), .B2(new_n666_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n728_), .A2(new_n574_), .A3(new_n263_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n735_), .B2(new_n339_), .ZN(new_n749_));
  XOR2_X1   g548(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n675_), .A2(new_n581_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT112), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n727_), .B2(new_n753_), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n679_), .A2(new_n619_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n726_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n513_), .B1(new_n756_), .B2(new_n440_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT113), .Z(new_n758_));
  NOR3_X1   g557(.A1(new_n619_), .A2(new_n652_), .A3(new_n642_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n695_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n440_), .A2(new_n513_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(G1336gat));
  INV_X1    g561(.A(new_n660_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n514_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n764_), .A2(new_n514_), .B1(new_n756_), .B2(new_n765_), .ZN(G1337gat));
  NOR3_X1   g565(.A1(new_n756_), .A2(new_n666_), .A3(new_n534_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n263_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G99gat), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g569(.A1(new_n756_), .A2(new_n339_), .A3(new_n535_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n660_), .A2(new_n440_), .A3(new_n339_), .A4(new_n263_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n421_), .A2(new_n423_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n411_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n370_), .B1(new_n436_), .B2(new_n402_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n390_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n660_), .A2(new_n430_), .B1(new_n777_), .B2(new_n339_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n778_), .B2(new_n263_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n690_), .B1(new_n779_), .B2(new_n565_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n691_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n675_), .B(new_n759_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(G106gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n771_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT115), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n788_), .B(new_n771_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n787_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1339gat));
  NAND2_X1  g592(.A1(new_n652_), .A2(new_n616_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n592_), .A2(KEYINPUT12), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n594_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n610_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n572_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(KEYINPUT118), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n611_), .B2(KEYINPUT55), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n611_), .A2(KEYINPUT55), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n608_), .A2(new_n573_), .A3(new_n610_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n571_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n571_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n794_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n477_), .A2(new_n478_), .A3(new_n482_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n474_), .A2(new_n478_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n489_), .B1(new_n485_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n490_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n616_), .B2(new_n612_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT57), .B(new_n649_), .C1(new_n810_), .C2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n649_), .B1(new_n810_), .B2(new_n816_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n493_), .A2(new_n614_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n571_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n571_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n816_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n649_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n614_), .A2(new_n815_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT58), .B(new_n830_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n565_), .A3(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n819_), .A2(new_n822_), .A3(new_n829_), .A4(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n643_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n733_), .B(new_n838_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n619_), .A2(new_n839_), .A3(KEYINPUT117), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT117), .B1(new_n619_), .B2(new_n839_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n688_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT54), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n688_), .B(new_n844_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n837_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT120), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n837_), .A2(new_n849_), .A3(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n666_), .A2(new_n444_), .A3(new_n440_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT121), .Z(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n652_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n847_), .A2(new_n858_), .A3(new_n853_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n493_), .B(new_n859_), .C1(new_n854_), .C2(KEYINPUT59), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(new_n856_), .ZN(G1340gat));
  NOR2_X1   g660(.A1(new_n619_), .A2(KEYINPUT60), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  MUX2_X1   g662(.A(KEYINPUT60), .B(new_n862_), .S(new_n863_), .Z(new_n864_));
  NAND3_X1  g663(.A1(new_n851_), .A2(new_n853_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n619_), .B(new_n859_), .C1(new_n854_), .C2(KEYINPUT59), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n863_), .B2(new_n868_), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n855_), .B2(new_n642_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n859_), .B1(new_n854_), .B2(KEYINPUT59), .ZN(new_n871_));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n642_), .B2(KEYINPUT123), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(KEYINPUT123), .B2(new_n872_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n870_), .B1(new_n871_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n855_), .B2(new_n650_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT124), .B(G134gat), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n688_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n871_), .B2(new_n878_), .ZN(G1343gat));
  NOR4_X1   g678(.A1(new_n763_), .A2(new_n263_), .A3(new_n440_), .A4(new_n339_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n851_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n652_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n620_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g684(.A1(new_n851_), .A2(new_n642_), .A3(new_n880_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n851_), .A2(new_n888_), .A3(new_n642_), .A4(new_n880_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n887_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n881_), .A2(new_n894_), .A3(new_n650_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n881_), .A2(new_n565_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n443_), .A2(new_n660_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n675_), .B(new_n900_), .C1(new_n837_), .C2(new_n846_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n652_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n902_), .A2(G169gat), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n903_), .A2(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(KEYINPUT62), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n904_), .B(new_n905_), .C1(new_n234_), .C2(new_n902_), .ZN(G1348gat));
  NOR3_X1   g705(.A1(new_n900_), .A2(new_n354_), .A3(new_n619_), .ZN(new_n907_));
  AOI21_X1  g706(.A(KEYINPUT126), .B1(new_n851_), .B2(new_n339_), .ZN(new_n908_));
  AOI221_X4 g707(.A(KEYINPUT120), .B1(new_n843_), .B2(new_n845_), .C1(new_n836_), .C2(new_n643_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n849_), .B1(new_n837_), .B2(new_n846_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT126), .B(new_n339_), .C1(new_n909_), .C2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n907_), .B1(new_n908_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT127), .ZN(new_n914_));
  AOI21_X1  g713(.A(G176gat), .B1(new_n901_), .B2(new_n620_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n913_), .A2(new_n914_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n907_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n339_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n918_), .B1(new_n921_), .B2(new_n911_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT127), .B1(new_n922_), .B2(new_n915_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n917_), .A2(new_n923_), .ZN(G1349gat));
  OAI211_X1 g723(.A(new_n642_), .B(new_n899_), .C1(new_n908_), .C2(new_n912_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n643_), .A2(new_n345_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n925_), .A2(new_n228_), .B1(new_n901_), .B2(new_n926_), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n901_), .A2(new_n202_), .A3(new_n650_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n901_), .A2(new_n565_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n229_), .ZN(G1351gat));
  INV_X1    g729(.A(new_n430_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n660_), .A2(new_n931_), .A3(new_n263_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n851_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n652_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g734(.A(new_n269_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n851_), .A2(new_n620_), .A3(new_n932_), .ZN(new_n937_));
  MUX2_X1   g736(.A(new_n936_), .B(G204gat), .S(new_n937_), .Z(G1353gat));
  NAND3_X1  g737(.A1(new_n851_), .A2(new_n642_), .A3(new_n932_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  AND2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n939_), .B2(new_n940_), .ZN(G1354gat));
  INV_X1    g742(.A(G218gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n933_), .A2(new_n944_), .A3(new_n650_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n933_), .A2(new_n565_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n947_), .B2(new_n944_), .ZN(G1355gat));
endmodule


