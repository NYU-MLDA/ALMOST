//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND4_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .A4(KEYINPUT65), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT65), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT7), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT8), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT10), .B(G99gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n206_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n214_), .A2(new_n215_), .A3(G85gat), .A4(G92gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n218_), .A2(new_n220_), .A3(new_n221_), .A4(new_n203_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G29gat), .B(G36gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT15), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G232gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT34), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT35), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n226_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n228_), .B(new_n233_), .C1(new_n223_), .C2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n231_), .A2(new_n232_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  XOR2_X1   g036(.A(G134gat), .B(G162gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G190gat), .B(G218gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT36), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n235_), .A2(new_n236_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n235_), .A2(new_n236_), .ZN(new_n246_));
  NOR4_X1   g045(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT36), .A4(new_n242_), .ZN(new_n247_));
  OR3_X1    g046(.A1(new_n244_), .A2(KEYINPUT37), .A3(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n243_), .B(KEYINPUT72), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n237_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT37), .B1(new_n250_), .B2(new_n247_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT73), .B(G15gat), .ZN(new_n253_));
  INV_X1    g052(.A(G22gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G1gat), .ZN(new_n256_));
  INV_X1    g055(.A(G8gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT14), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G8gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G71gat), .B(G78gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(KEYINPUT11), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT11), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n263_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G231gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G127gat), .B(G155gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT16), .ZN(new_n273_));
  INV_X1    g072(.A(G183gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G211gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT17), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n271_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT74), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT74), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT17), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n271_), .A2(new_n281_), .A3(new_n276_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n252_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT75), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n213_), .A2(new_n222_), .A3(new_n268_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G230gat), .A2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n268_), .B1(new_n213_), .B2(new_n222_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT68), .B1(new_n290_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n287_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n286_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(new_n291_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n288_), .B(KEYINPUT67), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT68), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n291_), .A2(new_n294_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G120gat), .B(G148gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(G204gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT5), .B(G176gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n305_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT13), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n313_), .A2(KEYINPUT69), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT69), .B1(new_n313_), .B2(new_n314_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT0), .ZN(new_n319_));
  INV_X1    g118(.A(G57gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT1), .ZN(new_n331_));
  INV_X1    g130(.A(G155gat), .ZN(new_n332_));
  INV_X1    g131(.A(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(new_n335_), .A3(new_n329_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G141gat), .ZN(new_n343_));
  INV_X1    g142(.A(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT3), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n349_), .A2(new_n350_), .B1(new_n338_), .B2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(KEYINPUT82), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n328_), .A2(new_n329_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n354_), .A2(KEYINPUT83), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT83), .B1(new_n354_), .B2(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n342_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G127gat), .B(G134gat), .Z(new_n359_));
  XOR2_X1   g158(.A(G113gat), .B(G120gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n361_), .B(new_n342_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT95), .A3(new_n364_), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n358_), .A2(KEYINPUT95), .A3(new_n362_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n325_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n358_), .A2(new_n325_), .A3(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT96), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT97), .B1(new_n367_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n365_), .A2(new_n366_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n369_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(KEYINPUT4), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT97), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n324_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n378_), .A2(new_n324_), .A3(new_n374_), .A4(new_n372_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  INV_X1    g182(.A(G190gat), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n274_), .A2(new_n384_), .A3(KEYINPUT23), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(G183gat), .B2(G190gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n383_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G169gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT22), .ZN(new_n392_));
  AOI21_X1  g191(.A(G176gat), .B1(new_n392_), .B2(KEYINPUT78), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G169gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(KEYINPUT78), .B2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(KEYINPUT79), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(KEYINPUT79), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n390_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT23), .B1(new_n274_), .B2(new_n384_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n385_), .B1(KEYINPUT77), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(KEYINPUT77), .B2(new_n400_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT25), .B(G183gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT26), .B(G190gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(G169gat), .B2(G176gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(G169gat), .B2(G176gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n399_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n385_), .A2(new_n387_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n389_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n398_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n383_), .B(new_n416_), .C1(new_n417_), .C2(new_n396_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT30), .B1(new_n418_), .B2(new_n410_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n413_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n412_), .B1(new_n399_), .B2(new_n411_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(new_n410_), .A3(KEYINPUT30), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G43gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT31), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n423_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n422_), .B1(new_n413_), .B2(new_n419_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n425_), .A2(new_n426_), .A3(new_n424_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n431_), .A2(new_n434_), .A3(KEYINPUT80), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n433_), .A3(new_n429_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n361_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT80), .B1(new_n431_), .B2(new_n434_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n362_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n382_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n446_), .B(KEYINPUT91), .Z(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(KEYINPUT19), .Z(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT92), .Z(new_n449_));
  XOR2_X1   g248(.A(G211gat), .B(G218gat), .Z(new_n450_));
  XOR2_X1   g249(.A(G197gat), .B(G204gat), .Z(new_n451_));
  INV_X1    g250(.A(KEYINPUT21), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n452_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT21), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n451_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G176gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n394_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n383_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n402_), .B2(new_n415_), .ZN(new_n463_));
  OAI22_X1  g262(.A1(new_n408_), .A2(KEYINPUT93), .B1(G169gat), .B2(G176gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(KEYINPUT93), .B2(new_n408_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n414_), .A2(new_n406_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n459_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT94), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n399_), .A2(new_n411_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n459_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n449_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G8gat), .B(G36gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT18), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G64gat), .ZN(new_n477_));
  INV_X1    g276(.A(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n471_), .B2(new_n472_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n463_), .A2(new_n467_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n448_), .B1(new_n482_), .B2(new_n459_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n474_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT27), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n469_), .A2(new_n449_), .A3(new_n473_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n448_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n455_), .A2(new_n451_), .A3(new_n457_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(new_n453_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n454_), .A2(new_n458_), .A3(KEYINPUT88), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(new_n482_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n489_), .B1(new_n481_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n480_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n487_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n469_), .A2(new_n473_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n449_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n484_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n479_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(new_n485_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n500_), .B1(KEYINPUT27), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G228gat), .A2(G233gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n358_), .A2(KEYINPUT29), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n494_), .B1(new_n512_), .B2(KEYINPUT87), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n358_), .A2(new_n514_), .A3(KEYINPUT29), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n517_));
  INV_X1    g316(.A(new_n341_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n330_), .A2(KEYINPUT1), .B1(new_n332_), .B2(new_n333_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n336_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n354_), .A2(new_n355_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT83), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n354_), .A2(KEYINPUT83), .A3(new_n355_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n520_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n517_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n358_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n528_));
  INV_X1    g327(.A(new_n511_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n472_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n510_), .B1(new_n516_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT87), .B1(new_n525_), .B2(new_n526_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n495_), .A3(new_n515_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n529_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n509_), .A3(new_n531_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(KEYINPUT85), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT89), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n525_), .A2(new_n526_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G22gat), .B(G50gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n533_), .A2(new_n545_), .A3(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n548_));
  INV_X1    g347(.A(new_n544_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n538_), .A3(KEYINPUT89), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n445_), .B(new_n508_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n538_), .A2(KEYINPUT89), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n546_), .A2(new_n544_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n550_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT90), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n507_), .B1(new_n560_), .B2(new_n551_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(KEYINPUT100), .A3(new_n445_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n368_), .A2(new_n369_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n324_), .B1(new_n376_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT98), .B1(new_n365_), .B2(new_n366_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n370_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT98), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n566_), .B(KEYINPUT99), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT99), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n570_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n323_), .B1(new_n367_), .B2(new_n564_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n375_), .A2(KEYINPUT33), .A3(new_n324_), .A4(new_n378_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n380_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .A4(new_n506_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n488_), .B2(new_n497_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n474_), .A2(new_n484_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(new_n581_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n444_), .B1(new_n563_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n382_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n560_), .B(new_n551_), .C1(new_n588_), .C2(new_n507_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n556_), .A2(new_n562_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n261_), .A2(new_n226_), .A3(new_n262_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT76), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT76), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n263_), .A2(new_n234_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n593_), .A2(new_n594_), .B1(new_n227_), .B2(new_n263_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n591_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n391_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G197gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n599_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR4_X1   g403(.A1(new_n285_), .A2(new_n317_), .A3(new_n590_), .A4(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n256_), .A3(new_n588_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT38), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n244_), .A2(new_n247_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT101), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n590_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n283_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n311_), .B(KEYINPUT13), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT69), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n603_), .A4(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n382_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n607_), .A2(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n605_), .A2(new_n257_), .A3(new_n507_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G8gat), .B1(new_n614_), .B2(new_n508_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT39), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(KEYINPUT39), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(G1325gat));
  INV_X1    g422(.A(new_n444_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G15gat), .B1(new_n614_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n605_), .A2(new_n627_), .A3(new_n444_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1326gat));
  OAI21_X1  g428(.A(G22gat), .B1(new_n614_), .B2(new_n563_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  INV_X1    g430(.A(new_n563_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n605_), .A2(new_n254_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1327gat));
  OAI211_X1 g433(.A(new_n283_), .B(new_n603_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n608_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n590_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G29gat), .B1(new_n637_), .B2(new_n588_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n252_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT43), .B1(new_n590_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n563_), .A2(new_n586_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n589_), .A3(new_n624_), .ZN(new_n642_));
  AND4_X1   g441(.A1(KEYINPUT100), .A2(new_n563_), .A3(new_n508_), .A4(new_n445_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT100), .B1(new_n561_), .B2(new_n445_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n252_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n635_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n650_), .A2(G29gat), .A3(new_n588_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n590_), .A2(KEYINPUT43), .A3(new_n639_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n646_), .B1(new_n645_), .B2(new_n252_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n638_), .B1(new_n651_), .B2(new_n656_), .ZN(G1328gat));
  AOI211_X1 g456(.A(new_n655_), .B(new_n635_), .C1(new_n640_), .C2(new_n647_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n508_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n637_), .A2(new_n663_), .A3(new_n507_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT45), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n661_), .A2(KEYINPUT102), .A3(new_n662_), .A4(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(KEYINPUT102), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n662_), .A2(KEYINPUT102), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n663_), .B1(new_n659_), .B2(new_n656_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n664_), .B(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n667_), .B(new_n668_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n666_), .A2(new_n672_), .ZN(G1329gat));
  NAND2_X1  g472(.A1(new_n637_), .A2(new_n444_), .ZN(new_n674_));
  INV_X1    g473(.A(G43gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n649_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n658_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n624_), .A2(new_n675_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT103), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  AND4_X1   g479(.A1(KEYINPUT103), .A2(new_n656_), .A3(new_n650_), .A4(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n676_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT47), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n676_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n637_), .B2(new_n632_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n632_), .A2(G50gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n678_), .B2(new_n688_), .ZN(G1331gat));
  NAND2_X1  g488(.A1(new_n317_), .A2(new_n604_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n285_), .A3(new_n590_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n320_), .A3(new_n588_), .ZN(new_n692_));
  NOR4_X1   g491(.A1(new_n690_), .A2(new_n609_), .A3(new_n590_), .A4(new_n283_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n588_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(new_n320_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n693_), .B2(new_n507_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT48), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n691_), .A2(new_n696_), .A3(new_n507_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n693_), .B2(new_n444_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n691_), .A2(new_n701_), .A3(new_n444_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n691_), .A2(new_n707_), .A3(new_n632_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n693_), .A2(new_n632_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G78gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT105), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n712_), .A3(G78gat), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n711_), .A2(KEYINPUT50), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT50), .B1(new_n711_), .B2(new_n713_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n708_), .B1(new_n714_), .B2(new_n715_), .ZN(G1335gat));
  NAND3_X1  g515(.A1(new_n317_), .A2(new_n283_), .A3(new_n604_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n717_), .A2(new_n636_), .A3(new_n590_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n588_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT106), .Z(new_n720_));
  INV_X1    g519(.A(new_n717_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n648_), .A2(KEYINPUT107), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT107), .B1(new_n648_), .B2(new_n721_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n382_), .A2(new_n322_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n720_), .B1(new_n724_), .B2(new_n725_), .ZN(G1336gat));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(G92gat), .A3(new_n507_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n718_), .A2(new_n507_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n478_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(KEYINPUT108), .A3(new_n478_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n727_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n728_), .A2(KEYINPUT109), .A3(new_n734_), .A4(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1337gat));
  NAND3_X1  g537(.A1(new_n718_), .A2(new_n219_), .A3(new_n444_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n648_), .A2(new_n444_), .A3(new_n721_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n205_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n648_), .A2(new_n632_), .A3(new_n721_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n648_), .A2(KEYINPUT110), .A3(new_n632_), .A4(new_n721_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n206_), .B1(new_n747_), .B2(KEYINPUT52), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n746_), .A3(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(KEYINPUT52), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n750_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n745_), .A2(new_n752_), .A3(new_n746_), .A4(new_n748_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n718_), .A2(new_n206_), .A3(new_n632_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT53), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n751_), .A2(new_n757_), .A3(new_n753_), .A4(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  NOR3_X1   g558(.A1(new_n252_), .A2(new_n283_), .A3(new_n603_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n612_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(new_n612_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n595_), .A2(new_n596_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n591_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n591_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n602_), .B1(new_n598_), .B2(new_n768_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n599_), .A2(new_n602_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n311_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n290_), .A2(new_n295_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n303_), .A2(new_n286_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n772_), .A2(KEYINPUT55), .B1(new_n297_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n296_), .A2(new_n775_), .A3(new_n304_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n310_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n296_), .A2(new_n775_), .A3(new_n304_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n773_), .A2(new_n297_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n300_), .A2(new_n303_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n775_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n310_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n777_), .A2(KEYINPUT112), .A3(KEYINPUT56), .A4(new_n310_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n305_), .A2(new_n310_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n603_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n771_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n765_), .B1(new_n793_), .B2(new_n608_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n310_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n786_), .B(new_n309_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(KEYINPUT112), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n791_), .B1(new_n797_), .B2(new_n780_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT57), .B(new_n636_), .C1(new_n798_), .C2(new_n771_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n790_), .A2(new_n770_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n787_), .B2(new_n778_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n252_), .B1(new_n801_), .B2(KEYINPUT58), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n790_), .A2(new_n770_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(KEYINPUT58), .C1(new_n796_), .C2(new_n795_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT113), .B1(new_n802_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n795_), .A2(new_n796_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n800_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n252_), .A4(new_n804_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n794_), .A2(new_n799_), .A3(new_n806_), .A4(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n764_), .B1(new_n812_), .B2(new_n283_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n561_), .A2(new_n588_), .A3(new_n444_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n603_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT59), .B1(new_n813_), .B2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n794_), .A2(new_n799_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n802_), .A2(new_n805_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n283_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n764_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n814_), .A2(KEYINPUT59), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n818_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT114), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n818_), .A2(new_n825_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n604_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n817_), .B1(new_n830_), .B2(new_n816_), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n826_), .B2(new_n613_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n815_), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n613_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(KEYINPUT60), .B2(new_n834_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n833_), .B2(new_n836_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT115), .B(new_n838_), .C1(new_n833_), .C2(new_n283_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n813_), .A2(new_n283_), .A3(new_n814_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(G127gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n827_), .A2(new_n829_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n283_), .A2(new_n838_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(G1342gat));
  AOI21_X1  g645(.A(G134gat), .B1(new_n815_), .B2(new_n609_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n252_), .A2(G134gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT116), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n844_), .B2(new_n849_), .ZN(G1343gat));
  XNOR2_X1  g649(.A(KEYINPUT118), .B(G141gat), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n812_), .A2(new_n283_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n822_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n563_), .A2(new_n444_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n507_), .A2(new_n382_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT117), .ZN(new_n858_));
  INV_X1    g657(.A(new_n855_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n813_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n856_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n852_), .B1(new_n863_), .B2(new_n603_), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n604_), .B(new_n851_), .C1(new_n858_), .C2(new_n862_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1344gat));
  XNOR2_X1  g665(.A(KEYINPUT119), .B(G148gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n863_), .B2(new_n317_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n613_), .B(new_n867_), .C1(new_n858_), .C2(new_n862_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1345gat));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT120), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n863_), .B2(new_n611_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  AOI211_X1 g674(.A(new_n283_), .B(new_n875_), .C1(new_n858_), .C2(new_n862_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1346gat));
  NAND3_X1  g676(.A1(new_n863_), .A2(new_n333_), .A3(new_n609_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n639_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n333_), .B2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g679(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n508_), .A2(new_n588_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n624_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n632_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n823_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT121), .B1(new_n887_), .B2(new_n604_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n391_), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n887_), .A2(KEYINPUT121), .A3(new_n604_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n881_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  OR3_X1    g691(.A1(new_n887_), .A2(KEYINPUT121), .A3(new_n604_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n881_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n893_), .A2(new_n888_), .A3(new_n889_), .A4(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n887_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n394_), .A3(new_n603_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n895_), .A3(new_n897_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n896_), .B2(new_n317_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n632_), .B1(new_n853_), .B2(new_n822_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n613_), .A2(new_n460_), .A3(new_n885_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n884_), .A2(new_n611_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n900_), .B2(new_n906_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n813_), .A2(KEYINPUT123), .A3(new_n632_), .A4(new_n905_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n907_), .A2(new_n908_), .A3(G183gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n887_), .A2(new_n404_), .A3(new_n283_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n903_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n910_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n813_), .A2(new_n632_), .A3(new_n905_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n274_), .B1(new_n913_), .B2(new_n904_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n912_), .B(KEYINPUT124), .C1(new_n908_), .C2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n915_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n887_), .B2(new_n639_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n609_), .A2(new_n405_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n887_), .B2(new_n918_), .ZN(G1351gat));
  NAND2_X1  g718(.A1(new_n860_), .A2(new_n882_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n603_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g722(.A1(new_n920_), .A2(new_n613_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(G204gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(G204gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT126), .Z(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OR3_X1    g728(.A1(new_n924_), .A2(new_n926_), .A3(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n924_), .B2(new_n926_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1353gat));
  NAND3_X1  g731(.A1(new_n860_), .A2(new_n611_), .A3(new_n882_), .ZN(new_n933_));
  OR2_X1    g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT63), .B(G211gat), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n860_), .A2(new_n611_), .A3(new_n882_), .A4(new_n937_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n935_), .A2(new_n936_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n936_), .B1(new_n935_), .B2(new_n938_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n920_), .B2(new_n639_), .ZN(new_n942_));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n609_), .A2(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n942_), .B1(new_n920_), .B2(new_n944_), .ZN(G1355gat));
endmodule


