//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT83), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT84), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT82), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  INV_X1    g011(.A(G176gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT24), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT80), .B(G183gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT25), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n218_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT81), .B1(new_n218_), .B2(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n221_), .A2(G183gat), .B1(new_n218_), .B2(G190gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n209_), .A2(new_n215_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(new_n203_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n204_), .A2(new_n207_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n213_), .B1(new_n230_), .B2(KEYINPUT85), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G169gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(G169gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT86), .B(G43gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT87), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G15gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n238_), .B(new_n241_), .Z(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT88), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(new_n244_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT31), .Z(new_n250_));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  OR2_X1    g051(.A1(new_n242_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT94), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(G204gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(G211gat), .B(G218gat), .Z(new_n261_));
  INV_X1    g060(.A(G204gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT95), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  OR4_X1    g062(.A1(new_n256_), .A2(new_n260_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(G197gat), .ZN(new_n265_));
  OAI221_X1 g064(.A(new_n265_), .B1(new_n262_), .B2(new_n259_), .C1(new_n261_), .C2(new_n256_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT95), .A2(KEYINPUT21), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n261_), .A2(new_n267_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G141gat), .ZN(new_n270_));
  INV_X1    g069(.A(G148gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT90), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n272_), .A2(KEYINPUT3), .B1(new_n274_), .B2(KEYINPUT2), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n273_), .B(KEYINPUT89), .ZN(new_n276_));
  OAI221_X1 g075(.A(new_n275_), .B1(KEYINPUT3), .B2(new_n272_), .C1(new_n276_), .C2(KEYINPUT2), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G155gat), .B(G162gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT91), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT1), .B2(new_n278_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n269_), .B1(new_n285_), .B2(KEYINPUT29), .ZN(new_n286_));
  INV_X1    g085(.A(G233gat), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(KEYINPUT93), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(KEYINPUT93), .ZN(new_n289_));
  OAI21_X1  g088(.A(G228gat), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n286_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G78gat), .B(G106gat), .Z(new_n292_));
  OR2_X1    g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n292_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n285_), .A2(KEYINPUT29), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT28), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G22gat), .B(G50gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n298_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n285_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(new_n249_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n306_), .B2(new_n245_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT4), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n306_), .A2(KEYINPUT4), .A3(new_n249_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT101), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n308_), .A2(new_n316_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G29gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G57gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  NAND3_X1  g123(.A1(new_n320_), .A2(KEYINPUT33), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT33), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n318_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n324_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n325_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G169gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n213_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n333_), .B(new_n335_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n210_), .A2(new_n224_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n215_), .A2(new_n228_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n269_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n344_), .B(KEYINPUT20), .C1(new_n343_), .C2(new_n235_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n336_), .A2(new_n269_), .A3(new_n341_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT97), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n351_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n343_), .B2(new_n235_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n349_), .B1(new_n356_), .B2(new_n348_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT99), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT98), .B(KEYINPUT18), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(KEYINPUT100), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n358_), .A2(new_n364_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT100), .B1(new_n357_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n332_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n320_), .A2(new_n324_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n329_), .A2(new_n330_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n350_), .A2(new_n355_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n348_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n345_), .B2(new_n375_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n357_), .B2(new_n378_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n373_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n305_), .B1(new_n370_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n304_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n302_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n369_), .A2(new_n385_), .A3(new_n365_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n385_), .B1(new_n377_), .B2(new_n367_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n366_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n384_), .A2(new_n373_), .A3(new_n386_), .A4(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n255_), .B1(new_n382_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n255_), .A2(new_n373_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n384_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G85gat), .ZN(new_n395_));
  INV_X1    g194(.A(G92gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G85gat), .A2(G92gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G99gat), .A2(G106gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G99gat), .A3(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT7), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n400_), .B1(new_n408_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT8), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT69), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n402_), .A2(new_n404_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n409_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n412_), .A2(new_n413_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT66), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423_));
  INV_X1    g222(.A(G99gat), .ZN(new_n424_));
  INV_X1    g223(.A(G106gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n411_), .A3(new_n410_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT66), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n419_), .A4(new_n409_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n399_), .A2(new_n417_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n414_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n435_), .B(KEYINPUT8), .C1(new_n436_), .C2(new_n400_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n427_), .A2(new_n419_), .A3(new_n409_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n430_), .B1(new_n438_), .B2(KEYINPUT66), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(KEYINPUT67), .A3(new_n429_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n418_), .A2(new_n434_), .A3(new_n437_), .A4(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G29gat), .B(G36gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G43gat), .B(G50gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT64), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n397_), .B1(new_n445_), .B2(KEYINPUT9), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n445_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT10), .B(G99gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n419_), .B1(new_n449_), .B2(G106gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n441_), .A2(new_n444_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G232gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT34), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT35), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n419_), .A2(KEYINPUT68), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n409_), .A3(new_n427_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n399_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n435_), .B1(new_n461_), .B2(KEYINPUT8), .ZN(new_n462_));
  AOI211_X1 g261(.A(KEYINPUT69), .B(new_n417_), .C1(new_n460_), .C2(new_n399_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND4_X1   g263(.A1(KEYINPUT67), .A2(new_n422_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT67), .B1(new_n439_), .B2(new_n429_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n451_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n444_), .B(KEYINPUT15), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n453_), .B(new_n457_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n455_), .A2(KEYINPUT35), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(KEYINPUT72), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n441_), .A2(new_n452_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n456_), .B1(new_n476_), .B2(new_n469_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n473_), .A3(new_n453_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G190gat), .B(G218gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT73), .ZN(new_n480_));
  XOR2_X1   g279(.A(G134gat), .B(G162gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT74), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI211_X1 g288(.A(new_n485_), .B(new_n487_), .C1(new_n475_), .C2(new_n478_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT103), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT103), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n497_));
  AND2_X1   g296(.A1(G230gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G64gat), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n499_), .A2(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n501_), .A2(new_n502_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n441_), .B2(new_n452_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT70), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508_));
  INV_X1    g307(.A(new_n505_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n508_), .B1(new_n476_), .B2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n498_), .B(new_n507_), .C1(new_n510_), .C2(new_n506_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n498_), .B1(new_n468_), .B2(new_n505_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n476_), .B2(new_n509_), .ZN(new_n514_));
  AOI211_X1 g313(.A(KEYINPUT12), .B(new_n505_), .C1(new_n441_), .C2(new_n452_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n512_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G120gat), .B(G148gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G176gat), .B(G204gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n511_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n511_), .B2(new_n516_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n497_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n511_), .A2(new_n516_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n521_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n511_), .A2(new_n516_), .A3(new_n522_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT13), .A3(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G8gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G15gat), .ZN(new_n535_));
  INV_X1    g334(.A(G22gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G15gat), .A2(G22gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G1gat), .A2(G8gat), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n537_), .A2(new_n538_), .B1(KEYINPUT14), .B2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n469_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n444_), .A3(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT78), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n544_), .A2(new_n545_), .A3(new_n549_), .A4(new_n546_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n543_), .B(new_n444_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n548_), .B(new_n550_), .C1(new_n546_), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT79), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G113gat), .B(G141gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n554_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n531_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n505_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(new_n543_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(G183gat), .B(G211gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n564_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n571_), .B2(new_n564_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n560_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n394_), .A2(new_n496_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G1gat), .B1(new_n577_), .B2(new_n373_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT38), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n390_), .A2(new_n393_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT102), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n471_), .A2(new_n474_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n473_), .B1(new_n477_), .B2(new_n453_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT74), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n584_), .A2(new_n487_), .B1(new_n585_), .B2(new_n483_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  INV_X1    g387(.A(new_n490_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n588_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n591_), .B(new_n592_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n530_), .A2(new_n590_), .A3(new_n593_), .A4(new_n574_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n580_), .A2(new_n581_), .A3(new_n558_), .A4(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n558_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT102), .B1(new_n597_), .B2(new_n594_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n373_), .A2(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n579_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n600_), .B2(new_n579_), .ZN(new_n603_));
  OAI221_X1 g402(.A(new_n578_), .B1(new_n579_), .B2(new_n600_), .C1(new_n602_), .C2(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n576_), .A2(KEYINPUT106), .A3(new_n391_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G8gat), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT106), .B1(new_n576_), .B2(new_n391_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n611_), .A2(KEYINPUT39), .A3(G8gat), .A4(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n391_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(G8gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n596_), .A2(new_n598_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT105), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n605_), .B1(new_n613_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n616_), .B(KEYINPUT105), .Z(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(KEYINPUT40), .A3(new_n612_), .A4(new_n610_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(G1325gat));
  AOI21_X1  g420(.A(new_n535_), .B1(new_n576_), .B2(new_n255_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n580_), .A2(new_n558_), .A3(new_n595_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n535_), .A3(new_n255_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(G1326gat));
  AOI21_X1  g426(.A(new_n536_), .B1(new_n576_), .B2(new_n384_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT42), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n536_), .A3(new_n384_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1327gat));
  NOR2_X1   g430(.A1(new_n491_), .A2(new_n574_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n580_), .A2(new_n558_), .A3(new_n530_), .A4(new_n632_), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n633_), .A2(G29gat), .A3(new_n373_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n590_), .A2(new_n593_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n574_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT43), .B(new_n635_), .C1(new_n390_), .C2(new_n393_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n560_), .A4(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n373_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n574_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(KEYINPUT44), .A3(new_n560_), .A4(new_n640_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT107), .ZN(new_n648_));
  OAI21_X1  g447(.A(G29gat), .B1(new_n647_), .B2(KEYINPUT107), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n634_), .B1(new_n648_), .B2(new_n649_), .ZN(G1328gat));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n391_), .A3(new_n646_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G36gat), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n614_), .A2(KEYINPUT108), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n386_), .A2(KEYINPUT108), .A3(new_n388_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(G36gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n633_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT45), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n652_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n659_), .A3(KEYINPUT46), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  NAND3_X1  g463(.A1(new_n643_), .A2(new_n255_), .A3(new_n646_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G43gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n255_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n633_), .A2(G43gat), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n666_), .A2(KEYINPUT47), .A3(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1330gat));
  NAND3_X1  g472(.A1(new_n643_), .A2(new_n384_), .A3(new_n646_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G50gat), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n305_), .A2(G50gat), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT109), .Z(new_n677_));
  OR2_X1    g476(.A1(new_n633_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n675_), .A2(KEYINPUT110), .A3(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1331gat));
  NOR3_X1   g482(.A1(new_n394_), .A2(new_n558_), .A3(new_n530_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n590_), .A2(new_n593_), .A3(new_n574_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n644_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G57gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n580_), .A2(new_n495_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n531_), .A2(new_n559_), .A3(new_n574_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n373_), .A2(new_n690_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n689_), .A2(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n655_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n686_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n693_), .A2(new_n697_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G64gat), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT48), .B(new_n696_), .C1(new_n693_), .C2(new_n697_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(new_n698_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n686_), .A2(new_n708_), .A3(new_n255_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n693_), .A2(new_n255_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G71gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n713_), .B2(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n686_), .A2(new_n716_), .A3(new_n384_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n693_), .A2(new_n384_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G78gat), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT50), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT50), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1335gat));
  AND2_X1   g521(.A1(new_n684_), .A2(new_n632_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n395_), .A3(new_n644_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n530_), .A2(new_n558_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n645_), .A2(new_n640_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n644_), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n724_), .B1(new_n730_), .B2(new_n395_), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n723_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n728_), .A2(new_n697_), .A3(new_n729_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n396_), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n726_), .B2(new_n667_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n449_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n723_), .A2(new_n255_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n723_), .A2(new_n425_), .A3(new_n384_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n645_), .A2(new_n384_), .A3(new_n640_), .A4(new_n725_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(G106gat), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n741_), .B2(G106gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n740_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n740_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  INV_X1    g549(.A(G113gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n685_), .A2(new_n752_), .A3(new_n559_), .A4(new_n530_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT54), .B1(new_n594_), .B2(new_n558_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n546_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n546_), .B2(new_n551_), .ZN(new_n757_));
  MUX2_X1   g556(.A(new_n757_), .B(new_n552_), .S(new_n557_), .Z(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n528_), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n514_), .A2(new_n515_), .B1(new_n476_), .B2(new_n509_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n498_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n516_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n512_), .B(KEYINPUT55), .C1(new_n514_), .C2(new_n515_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n521_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n521_), .ZN(new_n767_));
  OAI211_X1 g566(.A(KEYINPUT58), .B(new_n759_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n635_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n521_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n521_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT58), .B1(new_n774_), .B2(new_n759_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT116), .B1(new_n769_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n558_), .A2(new_n528_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n758_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n758_), .B(KEYINPUT115), .C1(new_n523_), .C2(new_n524_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n491_), .B1(new_n778_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n759_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n635_), .A4(new_n768_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT57), .B(new_n491_), .C1(new_n778_), .C2(new_n783_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n776_), .A2(new_n786_), .A3(new_n791_), .A4(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n755_), .B1(new_n793_), .B2(new_n639_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n614_), .A2(new_n305_), .A3(new_n644_), .A4(new_n255_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n751_), .B1(new_n797_), .B2(new_n559_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n799_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n795_), .A2(KEYINPUT59), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n781_), .A2(new_n782_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n558_), .B(new_n528_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n492_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n805_), .A2(KEYINPUT57), .B1(new_n775_), .B2(new_n769_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n806_), .A2(KEYINPUT118), .B1(KEYINPUT57), .B2(new_n805_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  OAI221_X1 g607(.A(new_n808_), .B1(new_n769_), .B2(new_n775_), .C1(new_n805_), .C2(KEYINPUT57), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n574_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n802_), .B1(new_n810_), .B2(new_n755_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT59), .B1(new_n794_), .B2(new_n795_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n559_), .A2(new_n751_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n800_), .A2(new_n801_), .B1(new_n813_), .B2(new_n814_), .ZN(G1340gat));
  NAND2_X1  g614(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n816_), .A2(new_n792_), .A3(new_n809_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n755_), .B1(new_n817_), .B2(new_n639_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n802_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n812_), .B(new_n531_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n811_), .A2(KEYINPUT119), .A3(new_n531_), .A4(new_n812_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(G120gat), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G120gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n530_), .A2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n796_), .B(new_n826_), .C1(G120gat), .C2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT120), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n796_), .B2(new_n574_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(G127gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n574_), .A2(KEYINPUT121), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(G127gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n813_), .B2(new_n838_), .ZN(G1342gat));
  NAND2_X1  g638(.A1(new_n813_), .A2(new_n635_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G134gat), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n495_), .A2(G134gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n797_), .B2(new_n842_), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n794_), .A2(new_n255_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(new_n644_), .A3(new_n384_), .A4(new_n655_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n559_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT122), .B(G141gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1344gat));
  NOR2_X1   g647(.A1(new_n845_), .A2(new_n530_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(new_n271_), .ZN(G1345gat));
  NOR2_X1   g649(.A1(new_n845_), .A2(new_n639_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n851_), .B(new_n852_), .Z(G1346gat));
  INV_X1    g652(.A(new_n635_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G162gat), .B1(new_n845_), .B2(new_n854_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n495_), .A2(G162gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n845_), .B2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n655_), .A2(new_n392_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n305_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n818_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n558_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n334_), .A3(new_n558_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT62), .B1(new_n862_), .B2(G169gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n858_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n862_), .A2(G169gat), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n870_), .A2(KEYINPUT123), .A3(new_n864_), .A4(new_n863_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n871_), .ZN(G1348gat));
  INV_X1    g671(.A(new_n861_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n213_), .B1(new_n873_), .B2(new_n530_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n794_), .A2(new_n384_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n859_), .A2(G176gat), .A3(new_n531_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n874_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n874_), .B(KEYINPUT124), .C1(new_n876_), .C2(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1349gat));
  NOR2_X1   g681(.A1(new_n639_), .A2(new_n337_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n875_), .A2(new_n574_), .A3(new_n859_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n861_), .A2(new_n883_), .B1(new_n884_), .B2(new_n216_), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n873_), .B2(new_n854_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n861_), .A2(new_n338_), .A3(new_n496_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1351gat));
  NOR3_X1   g687(.A1(new_n655_), .A2(new_n644_), .A3(new_n305_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n844_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n559_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT125), .B(G197gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1352gat));
  NOR2_X1   g692(.A1(new_n890_), .A2(new_n530_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n262_), .ZN(G1353gat));
  INV_X1    g694(.A(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n574_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  XOR2_X1   g700(.A(KEYINPUT126), .B(G218gat), .Z(new_n902_));
  NOR3_X1   g701(.A1(new_n890_), .A2(new_n854_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n896_), .A2(new_n496_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n902_), .ZN(G1355gat));
endmodule


