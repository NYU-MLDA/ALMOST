//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n209_), .A2(new_n211_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n217_), .A3(new_n216_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n207_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n215_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n204_), .A2(KEYINPUT9), .A3(new_n206_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n206_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT9), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n221_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT64), .B1(new_n230_), .B2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n209_), .A2(new_n211_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n229_), .A4(new_n228_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n225_), .A2(KEYINPUT66), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n225_), .B2(new_n239_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT67), .B(G71gat), .ZN(new_n245_));
  INV_X1    g044(.A(G78gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n246_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT68), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n252_), .A3(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n245_), .B(G78gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n256_), .A2(new_n244_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  OR3_X1    g057(.A1(new_n242_), .A2(KEYINPUT69), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G230gat), .ZN(new_n260_));
  INV_X1    g059(.A(G233gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n258_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n228_), .A2(new_n229_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n237_), .B1(new_n265_), .B2(new_n236_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n238_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n216_), .A2(new_n217_), .ZN(new_n269_));
  AOI211_X1 g068(.A(KEYINPUT8), .B(new_n268_), .C1(new_n269_), .C2(new_n221_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n223_), .B1(new_n222_), .B2(new_n207_), .ZN(new_n271_));
  OAI22_X1  g070(.A1(new_n266_), .A2(new_n267_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n225_), .A2(new_n239_), .A3(KEYINPUT66), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n258_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n276_), .A3(KEYINPUT69), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(new_n262_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT12), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n225_), .B2(new_n239_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n264_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n262_), .B1(new_n242_), .B2(new_n258_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G120gat), .B(G148gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n278_), .A2(new_n284_), .A3(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT13), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(KEYINPUT13), .A3(new_n293_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G141gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G169gat), .B(G197gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  XNOR2_X1  g108(.A(G29gat), .B(G36gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G43gat), .B(G50gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT75), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n309_), .A2(new_n312_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G229gat), .A3(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n312_), .B(KEYINPUT15), .ZN(new_n317_));
  INV_X1    g116(.A(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n309_), .A2(new_n312_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n302_), .B1(new_n316_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n322_), .A3(new_n302_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(KEYINPUT76), .A3(new_n325_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G127gat), .B(G134gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT79), .ZN(new_n332_));
  XOR2_X1   g131(.A(G113gat), .B(G120gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT80), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G71gat), .B(G99gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G43gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT31), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n335_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G15gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT30), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n339_), .B(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT23), .ZN(new_n350_));
  INV_X1    g149(.A(G169gat), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT24), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n348_), .B(new_n350_), .C1(new_n346_), .C2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT77), .B(G183gat), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT25), .ZN(new_n358_));
  OR2_X1    g157(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n350_), .B1(G190gat), .B2(new_n357_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT81), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n343_), .A2(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n339_), .A2(new_n342_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n339_), .A2(new_n342_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n367_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G211gat), .B(G218gat), .Z(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT87), .B(G197gat), .Z(new_n376_));
  INV_X1    g175(.A(G204gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT21), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(G197gat), .B2(G204gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n375_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(G204gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  INV_X1    g183(.A(G197gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(G204gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n381_), .B1(new_n387_), .B2(KEYINPUT21), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT21), .A3(new_n375_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n366_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT25), .B(G183gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n355_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n354_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n350_), .B1(G183gat), .B2(G190gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n364_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n393_), .B1(new_n400_), .B2(new_n390_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n392_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n361_), .A2(new_n365_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n390_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n391_), .A2(new_n399_), .A3(new_n397_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n409_));
  AND3_X1   g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n405_), .B1(new_n410_), .B2(new_n404_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n403_), .A2(new_n393_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n407_), .A2(new_n408_), .A3(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n392_), .A2(new_n401_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n418_), .B(new_n420_), .C1(new_n421_), .C2(new_n404_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(KEYINPUT27), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n404_), .B1(new_n392_), .B2(new_n401_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n420_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n416_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT93), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n430_), .B(KEYINPUT27), .C1(new_n422_), .C2(new_n426_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n423_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G141gat), .ZN(new_n433_));
  INV_X1    g232(.A(G148gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT3), .ZN(new_n436_));
  OR3_X1    g235(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G141gat), .A2(G148gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT2), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n436_), .A2(new_n437_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(G155gat), .A2(G162gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT83), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT1), .ZN(new_n448_));
  AOI211_X1 g247(.A(KEYINPUT82), .B(new_n444_), .C1(new_n443_), .C2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n448_), .B2(new_n443_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(KEYINPUT82), .A3(new_n448_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n450_), .A2(new_n438_), .A3(new_n435_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n335_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n334_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n458_));
  NAND3_X1  g257(.A1(new_n335_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(G85gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT0), .B(G57gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n454_), .A2(new_n456_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n461_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n461_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n467_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n476_));
  OR3_X1    g275(.A1(new_n453_), .A2(KEYINPUT29), .A3(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n453_), .B2(KEYINPUT29), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G22gat), .B(G50gat), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT89), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT89), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n486_), .A3(new_n483_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n391_), .B1(new_n453_), .B2(KEYINPUT29), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n246_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n488_), .A2(new_n246_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT85), .B(G228gat), .Z(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT86), .B(G233gat), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(G106gat), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n491_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(new_n489_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n485_), .B(new_n487_), .C1(new_n496_), .C2(new_n499_), .ZN(new_n500_));
  OR3_X1    g299(.A1(new_n487_), .A2(new_n499_), .A3(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n432_), .A2(new_n475_), .A3(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n500_), .A2(new_n501_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT33), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n474_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT33), .B(new_n467_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n457_), .A2(new_n461_), .A3(new_n459_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n468_), .C1(new_n461_), .C2(new_n469_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n427_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .A4(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n424_), .A2(new_n425_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n512_), .B2(new_n411_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n475_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n504_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n374_), .B1(new_n503_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n432_), .A2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT94), .B(new_n423_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n475_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n373_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n502_), .A3(new_n524_), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n299_), .B(new_n330_), .C1(new_n517_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n309_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n258_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G127gat), .B(G155gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT16), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n529_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n529_), .A2(new_n535_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G134gat), .B(G162gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n317_), .A2(new_n272_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n549_), .B2(KEYINPUT71), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n274_), .A2(new_n312_), .A3(new_n275_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n548_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n551_), .A2(KEYINPUT71), .A3(new_n548_), .A4(new_n547_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n544_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n542_), .B(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n555_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT74), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n554_), .A2(KEYINPUT74), .A3(new_n555_), .A4(new_n558_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT37), .ZN(new_n564_));
  INV_X1    g363(.A(new_n556_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n565_), .A2(KEYINPUT37), .A3(new_n559_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n526_), .A2(new_n539_), .A3(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n569_));
  AOI21_X1  g368(.A(G1gat), .B1(new_n569_), .B2(KEYINPUT96), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n475_), .A3(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(KEYINPUT96), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n563_), .B(KEYINPUT97), .Z(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n517_), .B2(new_n525_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n326_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n299_), .A2(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n575_), .A2(new_n539_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n304_), .B1(new_n578_), .B2(new_n475_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT98), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n573_), .A2(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(new_n521_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n568_), .A2(new_n305_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(G8gat), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n585_), .A2(KEYINPUT39), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(KEYINPUT39), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n583_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n588_), .B(new_n590_), .ZN(G1325gat));
  INV_X1    g390(.A(G15gat), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n578_), .B2(new_n373_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT41), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n568_), .A2(new_n592_), .A3(new_n373_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(G1326gat));
  INV_X1    g395(.A(G22gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n578_), .B2(new_n504_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT42), .Z(new_n599_));
  NAND3_X1  g398(.A1(new_n568_), .A2(new_n597_), .A3(new_n504_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(G1327gat));
  INV_X1    g400(.A(new_n563_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n539_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n526_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(G29gat), .B1(new_n605_), .B2(new_n475_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n567_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n511_), .A2(new_n515_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n502_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n502_), .A2(new_n475_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n429_), .A2(new_n431_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n423_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n373_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n504_), .B(new_n523_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT43), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n567_), .B1(new_n517_), .B2(new_n525_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n539_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n577_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT100), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT44), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n620_), .A2(KEYINPUT44), .A3(new_n623_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n475_), .A2(G29gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n606_), .B1(new_n628_), .B2(new_n629_), .ZN(G1328gat));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n582_), .A3(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G36gat), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n604_), .A2(G36gat), .A3(new_n521_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT45), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT46), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(KEYINPUT46), .A3(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1329gat));
  NAND4_X1  g439(.A1(new_n626_), .A2(G43gat), .A3(new_n373_), .A4(new_n627_), .ZN(new_n641_));
  INV_X1    g440(.A(G43gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n604_), .B2(new_n374_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g444(.A1(new_n604_), .A2(G50gat), .A3(new_n502_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n626_), .A2(new_n504_), .A3(new_n627_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n648_));
  OAI21_X1  g447(.A(G50gat), .B1(new_n647_), .B2(KEYINPUT101), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(G1331gat));
  AND3_X1   g449(.A1(new_n328_), .A2(new_n539_), .A3(new_n329_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n575_), .A2(new_n299_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n475_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n326_), .B1(new_n517_), .B2(new_n525_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n567_), .A2(new_n539_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT102), .B1(new_n655_), .B2(new_n298_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n655_), .A2(KEYINPUT102), .A3(new_n298_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n522_), .A2(G57gat), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n653_), .A2(G57gat), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT103), .ZN(G1332gat));
  INV_X1    g460(.A(G64gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n652_), .B2(new_n582_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n662_), .A3(new_n582_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1333gat));
  INV_X1    g466(.A(G71gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n668_), .A3(new_n373_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n652_), .A2(new_n373_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G71gat), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(KEYINPUT49), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(KEYINPUT49), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1334gat));
  AOI21_X1  g475(.A(new_n246_), .B1(new_n652_), .B2(new_n504_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT50), .Z(new_n678_));
  NAND3_X1  g477(.A1(new_n658_), .A2(new_n246_), .A3(new_n504_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1335gat));
  NOR3_X1   g479(.A1(new_n298_), .A2(new_n602_), .A3(new_n539_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n654_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n202_), .B1(new_n682_), .B2(new_n522_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT106), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n299_), .A2(new_n621_), .A3(new_n576_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n620_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n616_), .A2(new_n619_), .A3(KEYINPUT107), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n685_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n522_), .A2(new_n202_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n684_), .B1(new_n689_), .B2(new_n690_), .ZN(G1336gat));
  OAI21_X1  g490(.A(new_n203_), .B1(new_n682_), .B2(new_n521_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT108), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n521_), .A2(new_n203_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n689_), .B2(new_n694_), .ZN(G1337gat));
  NAND2_X1  g494(.A1(new_n687_), .A2(new_n688_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n685_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n373_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G99gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n682_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n700_), .A2(new_n373_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n699_), .A2(KEYINPUT109), .A3(KEYINPUT51), .A4(new_n701_), .ZN(new_n702_));
  OR2_X1    g501(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n703_));
  NAND2_X1  g502(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n214_), .B1(new_n689_), .B2(new_n373_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n701_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n703_), .B(new_n704_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n702_), .A2(new_n707_), .ZN(G1338gat));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n215_), .A3(new_n504_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n685_), .A2(new_n502_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n215_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n615_), .A2(KEYINPUT43), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n617_), .A2(new_n618_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n710_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT110), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n714_), .A2(new_n715_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n715_), .B1(new_n714_), .B2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n709_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n709_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1339gat));
  AND3_X1   g525(.A1(new_n651_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT54), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n567_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(new_n567_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n315_), .A2(new_n320_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n302_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n319_), .A2(new_n321_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n732_), .B(new_n733_), .C1(new_n320_), .C2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n325_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n293_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n282_), .A2(KEYINPUT55), .A3(new_n283_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n272_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n258_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n739_), .B(new_n276_), .C1(new_n740_), .C2(KEYINPUT12), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n262_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT55), .B1(new_n282_), .B2(new_n283_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n738_), .B(new_n742_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n739_), .B1(new_n740_), .B2(KEYINPUT12), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n276_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(KEYINPUT111), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n291_), .B1(new_n745_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT56), .B(new_n291_), .C1(new_n745_), .C2(new_n750_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n737_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n567_), .B1(new_n755_), .B2(KEYINPUT58), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n755_), .B2(KEYINPUT112), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n759_), .B(new_n737_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n326_), .A2(new_n293_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n294_), .A2(new_n736_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n602_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n762_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n754_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n749_), .A2(KEYINPUT111), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n284_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n738_), .A4(new_n742_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n291_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n769_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n764_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(KEYINPUT57), .A3(new_n602_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n761_), .A2(new_n768_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n731_), .B1(new_n778_), .B2(new_n621_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n582_), .A2(new_n522_), .A3(new_n504_), .A4(new_n374_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(G113gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n326_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT57), .B1(new_n776_), .B2(new_n602_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n767_), .B(new_n563_), .C1(new_n775_), .C2(new_n764_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n539_), .B1(new_n789_), .B2(new_n761_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT59), .B(new_n780_), .C1(new_n790_), .C2(new_n731_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n786_), .A2(KEYINPUT114), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT114), .B1(new_n786_), .B2(new_n791_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n330_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n784_), .B1(new_n794_), .B2(new_n783_), .ZN(G1340gat));
  NOR2_X1   g594(.A1(new_n298_), .A2(KEYINPUT60), .ZN(new_n796_));
  INV_X1    g595(.A(G120gat), .ZN(new_n797_));
  MUX2_X1   g596(.A(KEYINPUT60), .B(new_n796_), .S(new_n797_), .Z(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n782_), .A2(KEYINPUT115), .A3(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n298_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G120gat), .B1(new_n804_), .B2(KEYINPUT116), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n806_), .B(new_n298_), .C1(new_n786_), .C2(new_n791_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT117), .B(new_n803_), .C1(new_n805_), .C2(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1341gat));
  INV_X1    g611(.A(G127gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n782_), .A2(new_n813_), .A3(new_n539_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n792_), .A2(new_n793_), .A3(new_n621_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n813_), .ZN(G1342gat));
  AOI21_X1  g615(.A(G134gat), .B1(new_n782_), .B2(new_n574_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n792_), .A2(new_n793_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT118), .B(G134gat), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n607_), .A2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT119), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n817_), .B1(new_n818_), .B2(new_n821_), .ZN(G1343gat));
  INV_X1    g621(.A(new_n779_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n522_), .A2(new_n502_), .A3(new_n373_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n521_), .A3(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n576_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(new_n433_), .ZN(G1344gat));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n298_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(new_n434_), .ZN(G1345gat));
  NOR2_X1   g628(.A1(new_n825_), .A2(new_n621_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT61), .B(G155gat), .Z(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1346gat));
  INV_X1    g631(.A(G162gat), .ZN(new_n833_));
  INV_X1    g632(.A(new_n574_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n825_), .B2(new_n834_), .ZN(new_n835_));
  XOR2_X1   g634(.A(new_n835_), .B(KEYINPUT120), .Z(new_n836_));
  NOR2_X1   g635(.A1(new_n567_), .A2(new_n833_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT121), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n825_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(G1347gat));
  NOR2_X1   g639(.A1(new_n779_), .A2(new_n504_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n521_), .A2(new_n523_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n326_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G169gat), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n844_), .A2(KEYINPUT122), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(KEYINPUT122), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT62), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n844_), .A2(KEYINPUT122), .A3(new_n848_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT22), .B(G169gat), .Z(new_n850_));
  OR2_X1    g649(.A1(new_n843_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n849_), .A3(new_n851_), .ZN(G1348gat));
  NAND2_X1  g651(.A1(new_n841_), .A2(new_n842_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G176gat), .B1(new_n854_), .B2(new_n299_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n841_), .B(KEYINPUT123), .Z(new_n856_));
  NOR4_X1   g655(.A1(new_n521_), .A2(new_n352_), .A3(new_n523_), .A4(new_n298_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1349gat));
  NOR3_X1   g657(.A1(new_n853_), .A2(new_n394_), .A3(new_n621_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n539_), .A3(new_n842_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n357_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n853_), .B2(new_n567_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n574_), .A2(new_n355_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n853_), .B2(new_n864_), .ZN(G1351gat));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n610_), .A2(new_n374_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT124), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n521_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n779_), .B2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT125), .B(new_n869_), .C1(new_n790_), .C2(new_n731_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n326_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n299_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g676(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n873_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT126), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n873_), .A2(new_n882_), .A3(new_n878_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n880_), .A2(new_n881_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n881_), .B1(new_n880_), .B2(new_n883_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1354gat));
  NAND2_X1  g685(.A1(new_n873_), .A2(new_n574_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT127), .B(G218gat), .Z(new_n888_));
  NOR2_X1   g687(.A1(new_n567_), .A2(new_n888_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n887_), .A2(new_n888_), .B1(new_n873_), .B2(new_n889_), .ZN(G1355gat));
endmodule


