//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(G43gat), .ZN(new_n202_));
  INV_X1    g001(.A(G50gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G29gat), .B(G36gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n207_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(KEYINPUT15), .A3(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  INV_X1    g016(.A(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G1gat), .B(G8gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n211_), .A2(new_n222_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n211_), .B(new_n222_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(new_n227_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(KEYINPUT83), .B2(new_n228_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234_));
  INV_X1    g033(.A(G169gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G197gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n233_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240_));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241_));
  INV_X1    g040(.A(G113gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G113gat), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n243_), .A2(G120gat), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(G120gat), .B1(new_n243_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n240_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n245_), .ZN(new_n249_));
  INV_X1    g048(.A(G120gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n243_), .A2(G120gat), .A3(new_n245_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT87), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT30), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(KEYINPUT30), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  INV_X1    g059(.A(G190gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT23), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G183gat), .A3(G190gat), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT86), .B(KEYINPUT23), .C1(new_n260_), .C2(new_n261_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n259_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT22), .B(G169gat), .ZN(new_n272_));
  INV_X1    g071(.A(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT85), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n235_), .A2(new_n273_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n280_), .A2(KEYINPUT24), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n262_), .A2(KEYINPUT84), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n262_), .A2(KEYINPUT84), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n266_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n271_), .A2(new_n275_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n257_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n255_), .A2(new_n288_), .A3(new_n256_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G43gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT31), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G71gat), .B(G99gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n294_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n301_));
  OR3_X1    g100(.A1(new_n295_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT96), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306_));
  INV_X1    g105(.A(G204gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT91), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT91), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G204gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT21), .B(new_n306_), .C1(new_n311_), .C2(G197gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(G211gat), .B(G218gat), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n311_), .B2(G197gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n312_), .B(new_n314_), .C1(new_n316_), .C2(KEYINPUT21), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(KEYINPUT21), .A3(new_n313_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n288_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n284_), .A2(KEYINPUT93), .A3(new_n268_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n322_));
  INV_X1    g121(.A(new_n268_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(new_n283_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n259_), .B1(new_n287_), .B2(new_n270_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n321_), .A2(new_n324_), .B1(new_n325_), .B2(new_n274_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n320_), .B(KEYINPUT20), .C1(new_n326_), .C2(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n319_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n317_), .A2(new_n318_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n289_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n329_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n331_), .A2(new_n333_), .A3(KEYINPUT20), .A4(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G8gat), .B(G36gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n305_), .B1(new_n336_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n325_), .A2(new_n274_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n284_), .A2(new_n268_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n345_), .A2(new_n319_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n319_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n329_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n329_), .B2(new_n327_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n344_), .B1(new_n350_), .B2(new_n342_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n330_), .A2(new_n335_), .A3(KEYINPUT96), .A4(new_n341_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n343_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT89), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT2), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(KEYINPUT89), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT88), .ZN(new_n359_));
  OAI22_X1  g158(.A1(new_n359_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  INV_X1    g160(.A(G141gat), .ZN(new_n362_));
  INV_X1    g161(.A(G148gat), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .A4(KEYINPUT88), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .A4(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n366_), .A2(KEYINPUT1), .B1(new_n362_), .B2(new_n363_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n354_), .A3(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n369_), .A2(new_n373_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n376_), .B1(new_n381_), .B2(KEYINPUT29), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G78gat), .B(G106gat), .Z(new_n386_));
  OAI22_X1  g185(.A1(new_n384_), .A2(new_n385_), .B1(KEYINPUT92), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n332_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G228gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n385_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n386_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n383_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n391_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT95), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n248_), .A2(new_n253_), .A3(new_n381_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n374_), .A2(new_n252_), .A3(new_n251_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n400_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n400_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n407_), .A3(new_n404_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G85gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(G1gat), .B(G29gat), .Z(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n406_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n330_), .A2(new_n335_), .A3(new_n341_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n341_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n344_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n353_), .A2(new_n398_), .A3(new_n416_), .A4(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n415_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n387_), .A2(new_n394_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n390_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n406_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n426_));
  AND4_X1   g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .A4(new_n395_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n427_), .A2(KEYINPUT97), .A3(new_n419_), .A4(new_n353_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n422_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n426_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n350_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n432_), .C1(new_n431_), .C2(new_n336_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n414_), .A2(KEYINPUT33), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n417_), .A2(new_n418_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n407_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n401_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n412_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n426_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .A4(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n398_), .B1(new_n433_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n304_), .B1(new_n429_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n304_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n398_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n353_), .A2(new_n419_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n444_), .A2(new_n416_), .A3(new_n445_), .A4(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n239_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT98), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G230gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT68), .B(G71gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G78gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(G57gat), .B(G64gat), .Z(new_n454_));
  INV_X1    g253(.A(KEYINPUT11), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n455_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G78gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n452_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n456_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  INV_X1    g265(.A(G92gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT64), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT9), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n465_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n473_), .B2(new_n469_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT65), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(KEYINPUT64), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n473_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT9), .B1(new_n465_), .B2(KEYINPUT64), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT65), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n482_), .A4(KEYINPUT66), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  OAI22_X1  g294(.A1(new_n495_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n494_), .A2(new_n496_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n468_), .A2(new_n473_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n491_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n497_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n489_), .B(new_n490_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n498_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n497_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n490_), .B1(new_n506_), .B2(new_n489_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n464_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT69), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n500_), .A2(new_n499_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n487_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT10), .B(G99gat), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n478_), .B(new_n479_), .C1(new_n513_), .C2(G106gat), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT67), .B1(new_n510_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n501_), .A3(new_n463_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n451_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n489_), .B(new_n522_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n506_), .B2(new_n489_), .ZN(new_n525_));
  OAI211_X1 g324(.A(KEYINPUT12), .B(new_n463_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n521_), .A2(new_n450_), .A3(new_n526_), .A4(new_n508_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n516_), .A2(new_n501_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n451_), .B1(new_n530_), .B2(new_n464_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n531_), .A2(new_n521_), .A3(KEYINPUT71), .A4(new_n526_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n519_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G148gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT73), .B(G120gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  OR2_X1    g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n449_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n222_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n463_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT17), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT81), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n548_), .B(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(KEYINPUT17), .B2(new_n553_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT82), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT70), .B1(new_n510_), .B2(new_n515_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n523_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n211_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n215_), .A2(new_n561_), .B1(new_n530_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n215_), .A2(new_n561_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n530_), .A2(new_n562_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT75), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT34), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT34), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n563_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G232gat), .ZN(new_n574_));
  INV_X1    g373(.A(G233gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n571_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n577_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n566_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n573_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n576_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(KEYINPUT35), .A3(new_n578_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G134gat), .ZN(new_n586_));
  INV_X1    g385(.A(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT77), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(new_n584_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT78), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT78), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n581_), .A2(new_n584_), .A3(new_n594_), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n581_), .A2(new_n584_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT79), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n588_), .B(KEYINPUT36), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n581_), .A2(new_n584_), .A3(KEYINPUT79), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n596_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n597_), .A2(new_n601_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n596_), .A2(KEYINPUT37), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n545_), .A2(new_n559_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n217_), .A3(new_n430_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT38), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n559_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(new_n604_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n544_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n239_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n416_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(G1324gat));
  OAI21_X1  g418(.A(G8gat), .B1(new_n617_), .B2(new_n446_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT39), .ZN(new_n621_));
  INV_X1    g420(.A(new_n446_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n610_), .A2(new_n218_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n617_), .B2(new_n304_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT41), .Z(new_n627_));
  INV_X1    g426(.A(new_n610_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n304_), .A2(G15gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(G1326gat));
  OAI21_X1  g429(.A(G22gat), .B1(new_n617_), .B2(new_n445_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT42), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n445_), .A2(G22gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n628_), .B2(new_n633_), .ZN(G1327gat));
  NOR3_X1   g433(.A1(new_n545_), .A2(new_n558_), .A3(new_n604_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G29gat), .B1(new_n635_), .B2(new_n430_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n443_), .A2(new_n447_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT37), .B1(new_n596_), .B2(new_n603_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n600_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n605_), .B(new_n639_), .C1(new_n593_), .C2(new_n595_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT43), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n637_), .B(new_n643_), .C1(new_n638_), .C2(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n616_), .A3(new_n559_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT99), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n558_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n650_), .A2(new_n651_), .A3(new_n616_), .A4(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n416_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n636_), .B1(new_n655_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n649_), .A2(new_n654_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n622_), .ZN(new_n660_));
  AOI211_X1 g459(.A(KEYINPUT101), .B(new_n446_), .C1(new_n649_), .C2(new_n654_), .ZN(new_n661_));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n635_), .A2(new_n662_), .A3(new_n622_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n657_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n660_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n659_), .A2(new_n658_), .A3(new_n622_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(G36gat), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n664_), .B(KEYINPUT45), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n671_), .A3(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(new_n672_), .ZN(G1329gat));
  INV_X1    g472(.A(G43gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n674_), .B(new_n304_), .C1(new_n649_), .C2(new_n654_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G43gat), .B1(new_n635_), .B2(new_n444_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n659_), .A2(G43gat), .A3(new_n444_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n635_), .A2(new_n444_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n674_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n677_), .A2(KEYINPUT47), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT47), .B1(new_n677_), .B2(new_n682_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n635_), .B2(new_n398_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n203_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n398_), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n544_), .A2(new_n238_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n613_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n638_), .A2(new_n640_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n416_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n614_), .A2(new_n689_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n416_), .B2(KEYINPUT103), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(KEYINPUT103), .B2(G57gat), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n693_), .A2(G57gat), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT104), .Z(G1332gat));
  OAI21_X1  g497(.A(G64gat), .B1(new_n694_), .B2(new_n446_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT105), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT48), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n692_), .A2(G64gat), .A3(new_n446_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n694_), .B2(new_n304_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT49), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n692_), .A2(G71gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n304_), .B2(new_n706_), .ZN(G1334gat));
  OAI21_X1  g506(.A(G78gat), .B1(new_n694_), .B2(new_n445_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT50), .Z(new_n709_));
  NOR3_X1   g508(.A1(new_n692_), .A2(G78gat), .A3(new_n445_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  AND2_X1   g510(.A1(new_n650_), .A2(new_n689_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(G85gat), .A3(new_n430_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n604_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(new_n637_), .A3(new_n559_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n689_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n466_), .B1(new_n716_), .B2(new_n416_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n713_), .A2(new_n717_), .ZN(G1336gat));
  NAND3_X1  g517(.A1(new_n712_), .A2(G92gat), .A3(new_n622_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n467_), .B1(new_n716_), .B2(new_n446_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT106), .ZN(G1337gat));
  NAND4_X1  g521(.A1(new_n715_), .A2(new_n481_), .A3(new_n444_), .A4(new_n689_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n712_), .A2(new_n444_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G99gat), .ZN(new_n726_));
  AOI211_X1 g525(.A(KEYINPUT107), .B(new_n493_), .C1(new_n712_), .C2(new_n444_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g528(.A1(new_n715_), .A2(new_n482_), .A3(new_n398_), .A4(new_n689_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n712_), .A2(new_n398_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G106gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT52), .B(new_n482_), .C1(new_n712_), .C2(new_n398_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g535(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n533_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n521_), .A2(new_n526_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n451_), .B1(new_n509_), .B2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n531_), .A2(new_n521_), .A3(KEYINPUT55), .A4(new_n526_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n533_), .A2(KEYINPUT109), .A3(new_n738_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  INV_X1    g549(.A(new_n540_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n741_), .A2(KEYINPUT110), .A3(new_n745_), .A4(new_n746_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .A4(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n542_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n225_), .A2(KEYINPUT112), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n223_), .A2(new_n756_), .A3(new_n224_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n227_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n237_), .B1(new_n230_), .B2(new_n226_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT113), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n228_), .A2(KEYINPUT83), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n237_), .C1(new_n228_), .C2(new_n231_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n764_), .A3(new_n759_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n763_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n749_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(KEYINPUT56), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT58), .B1(new_n754_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT116), .B1(new_n771_), .B2(new_n691_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n754_), .A2(new_n770_), .A3(KEYINPUT58), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT109), .B1(new_n533_), .B2(new_n738_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n740_), .B(new_n737_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n743_), .A2(new_n744_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n774_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n751_), .B1(new_n777_), .B2(KEYINPUT110), .ZN(new_n778_));
  INV_X1    g577(.A(new_n752_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n766_), .B(KEYINPUT114), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n780_), .A2(new_n542_), .A3(new_n781_), .A4(new_n753_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n609_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n772_), .A2(new_n773_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n781_), .A2(new_n543_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n238_), .A2(new_n542_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n794_), .B2(new_n750_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n793_), .B(KEYINPUT56), .C1(new_n778_), .C2(new_n779_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n791_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n789_), .B1(new_n797_), .B2(new_n714_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n792_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n540_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT111), .B1(new_n800_), .B2(new_n752_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n796_), .B(new_n799_), .C1(KEYINPUT56), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n790_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n789_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n604_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n559_), .B1(new_n787_), .B2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n691_), .A2(new_n544_), .A3(new_n239_), .A4(new_n558_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT54), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n622_), .A2(new_n416_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n304_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n810_), .A2(new_n445_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814_), .B2(new_n238_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n445_), .A3(new_n813_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n398_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT59), .A3(new_n813_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n239_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n815_), .B1(new_n821_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g621(.A(new_n250_), .B1(new_n544_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n814_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n250_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n544_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n250_), .ZN(G1341gat));
  AOI21_X1  g625(.A(G127gat), .B1(new_n814_), .B2(new_n558_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n820_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n558_), .A2(G127gat), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT117), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n827_), .B1(new_n828_), .B2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n814_), .B2(new_n714_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n691_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g633(.A1(new_n812_), .A2(new_n444_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n810_), .A2(new_n398_), .A3(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n239_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(new_n362_), .ZN(G1344gat));
  NOR2_X1   g637(.A1(new_n836_), .A2(new_n544_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT118), .B(G148gat), .Z(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1345gat));
  NOR2_X1   g640(.A1(new_n836_), .A2(new_n559_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT61), .B(G155gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  NOR3_X1   g643(.A1(new_n836_), .A2(new_n587_), .A3(new_n691_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n587_), .B1(new_n836_), .B2(new_n604_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT119), .B(new_n587_), .C1(new_n836_), .C2(new_n604_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n848_), .B2(new_n849_), .ZN(G1347gat));
  NOR3_X1   g649(.A1(new_n304_), .A2(new_n430_), .A3(new_n446_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n819_), .A2(new_n238_), .A3(new_n272_), .A4(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n238_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n810_), .A2(new_n445_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(G169gat), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n856_), .B2(G169gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n852_), .B1(new_n859_), .B2(new_n860_), .ZN(G1348gat));
  NAND3_X1  g660(.A1(new_n810_), .A2(new_n445_), .A3(new_n851_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n544_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT121), .B(G176gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1349gat));
  OAI211_X1 g664(.A(KEYINPUT122), .B(new_n260_), .C1(new_n862_), .C2(new_n559_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n278_), .B1(KEYINPUT122), .B2(new_n277_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n819_), .A2(new_n558_), .A3(new_n851_), .A4(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1350gat));
  OAI21_X1  g668(.A(G190gat), .B1(new_n862_), .B2(new_n691_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n714_), .A2(new_n276_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n862_), .B2(new_n871_), .ZN(G1351gat));
  NOR2_X1   g671(.A1(new_n444_), .A2(new_n446_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n804_), .B1(new_n803_), .B2(new_n604_), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n714_), .B(new_n789_), .C1(new_n802_), .C2(new_n790_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n772_), .A2(new_n786_), .A3(new_n773_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n558_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n809_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n427_), .B(new_n873_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n239_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(G197gat), .Z(G1352gat));
  NAND2_X1  g681(.A1(KEYINPUT123), .A2(G204gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n880_), .B2(new_n544_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  INV_X1    g684(.A(new_n427_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n308_), .B1(new_n310_), .B2(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n887_), .A2(new_n615_), .A3(new_n873_), .A4(new_n889_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n884_), .A2(new_n885_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n885_), .B1(new_n884_), .B2(new_n890_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1353gat));
  OR2_X1    g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT63), .B(G211gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n880_), .A2(new_n559_), .ZN(new_n896_));
  MUX2_X1   g695(.A(new_n894_), .B(new_n895_), .S(new_n896_), .Z(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n880_), .B2(new_n604_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n691_), .A2(new_n898_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT125), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n887_), .A2(new_n873_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT126), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n899_), .A2(new_n905_), .A3(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1355gat));
endmodule


