//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT78), .B(G8gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G1gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT14), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G1gat), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G50gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT73), .ZN(new_n211_));
  INV_X1    g010(.A(G43gat), .ZN(new_n212_));
  INV_X1    g011(.A(G29gat), .ZN(new_n213_));
  INV_X1    g012(.A(G36gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n211_), .A2(new_n212_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n212_), .B1(new_n211_), .B2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n209_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G43gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n211_), .A2(new_n212_), .A3(new_n218_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(G50gat), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n221_), .A2(new_n225_), .A3(KEYINPUT15), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n208_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT81), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n206_), .B(G8gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n226_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n208_), .A2(new_n237_), .A3(new_n230_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n208_), .A2(new_n226_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n233_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245_));
  INV_X1    g044(.A(G169gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G197gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT82), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT83), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n244_), .A2(new_n249_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n253_), .B2(KEYINPUT83), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n256_));
  INV_X1    g055(.A(G141gat), .ZN(new_n257_));
  INV_X1    g056(.A(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT3), .ZN(new_n260_));
  NAND3_X1  g059(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n256_), .A2(new_n262_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT29), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n267_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n272_), .B2(new_n267_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  OR3_X1    g076(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n278_), .A2(new_n279_), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n270_), .B(new_n271_), .C1(new_n277_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT28), .ZN(new_n283_));
  INV_X1    g082(.A(G22gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(G155gat), .B2(G162gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT88), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n276_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n272_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n291_), .A2(new_n280_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n271_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n283_), .A2(new_n284_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n284_), .B1(new_n283_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n209_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n282_), .A2(KEYINPUT28), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n292_), .B2(new_n271_), .ZN(new_n299_));
  OAI21_X1  g098(.A(G22gat), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n283_), .A2(new_n284_), .A3(new_n294_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(G50gat), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G78gat), .B(G106gat), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n270_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT29), .ZN(new_n308_));
  INV_X1    g107(.A(G204gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G197gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n248_), .A2(G204gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n314_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n315_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT90), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT90), .B1(new_n318_), .B2(new_n319_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n306_), .B1(new_n308_), .B2(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n322_), .B(new_n306_), .C1(new_n292_), .C2(new_n271_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n305_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n306_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n291_), .A2(new_n280_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n271_), .B1(new_n328_), .B2(new_n270_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n321_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT90), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n318_), .A2(new_n319_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n330_), .A2(new_n331_), .B1(new_n316_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n327_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n324_), .A3(new_n304_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n326_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT93), .B1(new_n303_), .B2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n326_), .A2(new_n335_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT93), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n302_), .A4(new_n297_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n324_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT91), .B1(new_n343_), .B2(new_n305_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n335_), .A2(new_n344_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT91), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n335_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n342_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n326_), .A2(new_n346_), .A3(new_n335_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n303_), .A2(new_n347_), .A3(new_n349_), .A4(new_n342_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n341_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(KEYINPUT84), .A3(new_n355_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT85), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT23), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(G183gat), .B2(G190gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n360_), .A2(new_n362_), .A3(new_n369_), .A4(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT26), .B(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n246_), .A2(new_n355_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT24), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(KEYINPUT24), .A3(new_n363_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n374_), .A2(new_n367_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n371_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n354_), .B1(new_n379_), .B2(new_n322_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT19), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n368_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n333_), .A2(new_n378_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n371_), .A2(new_n333_), .A3(new_n378_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n378_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n322_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(KEYINPUT20), .A3(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n382_), .B(KEYINPUT94), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  NAND3_X1  g196(.A1(new_n386_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n353_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n383_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n390_), .A2(new_n391_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT27), .B(new_n398_), .C1(new_n404_), .C2(new_n397_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n352_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G120gat), .ZN(new_n408_));
  OR2_X1    g207(.A1(G127gat), .A2(G134gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G127gat), .A2(G134gat), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(G127gat), .A2(G134gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G127gat), .A2(G134gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT86), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(G113gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n412_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n408_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT86), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n410_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n421_));
  OAI21_X1  g220(.A(G113gat), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n412_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(G120gat), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n328_), .A2(new_n427_), .A3(new_n270_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n328_), .B2(new_n270_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n292_), .A2(new_n427_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(KEYINPUT4), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT4), .B1(new_n328_), .B2(new_n270_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n434_), .A2(new_n425_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n434_), .B2(new_n425_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n433_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n430_), .A2(new_n439_), .A3(new_n432_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT98), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n433_), .A2(new_n438_), .A3(KEYINPUT98), .A4(new_n440_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G85gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT100), .B(G57gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n444_), .A2(new_n454_), .A3(new_n445_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n379_), .B(new_n425_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G15gat), .B(G43gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT31), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n458_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G71gat), .B(G99gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT30), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n461_), .B(new_n465_), .Z(new_n466_));
  NAND3_X1  g265(.A1(new_n407_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n455_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n307_), .A2(KEYINPUT96), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n292_), .A2(new_n427_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n425_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT102), .B1(new_n472_), .B2(new_n431_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT102), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n430_), .A2(new_n474_), .A3(new_n432_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n475_), .A3(new_n440_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n433_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n452_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n386_), .A2(new_n392_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n397_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n478_), .A2(new_n398_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n468_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n444_), .A2(new_n454_), .A3(new_n445_), .A4(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n469_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n397_), .A2(KEYINPUT32), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n404_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n386_), .A2(new_n392_), .A3(new_n486_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n444_), .A2(new_n454_), .A3(new_n445_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n454_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n487_), .B(new_n488_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n303_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT92), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n494_), .A2(new_n350_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n406_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n457_), .A2(new_n352_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n466_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT104), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n352_), .B1(new_n485_), .B2(new_n491_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n495_), .A2(new_n456_), .A3(new_n406_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT104), .B(new_n500_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n467_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G230gat), .A2(G233gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT11), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT65), .B(G71gat), .ZN(new_n510_));
  INV_X1    g309(.A(G78gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT65), .B(G71gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(G78gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT11), .A3(new_n512_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(KEYINPUT11), .A3(new_n512_), .A4(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n526_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT8), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n535_), .B(new_n526_), .C1(new_n529_), .C2(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n530_), .B(KEYINPUT6), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n524_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n526_), .A2(KEYINPUT9), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT10), .B(G99gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT64), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n542_), .B(new_n543_), .C1(new_n545_), .C2(G106gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n537_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT66), .B1(new_n523_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT64), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n544_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(G106gat), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n541_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n552_), .A2(new_n543_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT66), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n520_), .A2(new_n522_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(KEYINPUT67), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n523_), .A2(new_n547_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT67), .B1(new_n548_), .B2(new_n556_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n508_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT68), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n523_), .A2(KEYINPUT12), .A3(new_n547_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n553_), .A2(new_n555_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .A4(new_n507_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n563_), .A2(new_n565_), .A3(new_n568_), .A4(new_n507_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT69), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT68), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n573_), .B(new_n508_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n562_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G176gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n309_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n562_), .A2(new_n572_), .A3(new_n574_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT70), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n580_), .A2(new_n582_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n523_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n208_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n594_), .A2(new_n595_), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(KEYINPUT17), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n229_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT15), .B1(new_n221_), .B2(new_n225_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n547_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT74), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT74), .B(new_n547_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n610_), .A2(new_n611_), .B1(new_n235_), .B2(new_n553_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT71), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT35), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT75), .B1(new_n610_), .B2(new_n611_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(KEYINPUT35), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT72), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n612_), .B(new_n616_), .C1(new_n617_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n235_), .A2(new_n553_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n611_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT74), .B1(new_n230_), .B2(new_n547_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n616_), .B(new_n622_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT75), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n627_), .A3(new_n619_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n628_), .A3(KEYINPUT77), .ZN(new_n629_));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT76), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(G134gat), .ZN(new_n632_));
  INV_X1    g431(.A(G162gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(KEYINPUT36), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n621_), .A2(new_n628_), .A3(KEYINPUT77), .A4(new_n636_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n621_), .A2(new_n628_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT36), .A3(new_n635_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n640_), .A2(KEYINPUT37), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT37), .B1(new_n640_), .B2(new_n642_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n590_), .B(new_n605_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT80), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT80), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n255_), .B(new_n506_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT105), .ZN(new_n649_));
  INV_X1    g448(.A(G1gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n456_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n589_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n580_), .A2(new_n582_), .B1(KEYINPUT70), .B2(new_n584_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n255_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n590_), .A2(KEYINPUT106), .A3(new_n255_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n467_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n665_), .B2(new_n504_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n640_), .A2(new_n642_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n604_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n661_), .A2(new_n666_), .A3(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT107), .Z(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(new_n456_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n653_), .B(new_n654_), .C1(new_n650_), .C2(new_n672_), .ZN(G1324gat));
  INV_X1    g472(.A(new_n203_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n649_), .A2(new_n674_), .A3(new_n406_), .ZN(new_n675_));
  NOR4_X1   g474(.A1(new_n661_), .A2(new_n666_), .A3(new_n669_), .A4(new_n497_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n676_), .A2(KEYINPUT108), .A3(new_n207_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT108), .B1(new_n676_), .B2(new_n207_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n675_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n675_), .B(KEYINPUT40), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1325gat));
  OR3_X1    g485(.A1(new_n648_), .A2(G15gat), .A3(new_n500_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(new_n466_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n688_), .B2(G15gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(G1326gat));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n671_), .A2(new_n352_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G22gat), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT42), .B(new_n284_), .C1(new_n671_), .C2(new_n352_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n352_), .A2(new_n284_), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n694_), .A2(new_n695_), .B1(new_n648_), .B2(new_n696_), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n667_), .A2(new_n604_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n700_), .A2(new_n666_), .A3(new_n657_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n213_), .A3(new_n456_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n659_), .A2(new_n604_), .A3(new_n660_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT37), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n667_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n640_), .A2(KEYINPUT37), .A3(new_n642_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n705_), .B1(new_n506_), .B2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n666_), .A2(KEYINPUT43), .A3(new_n709_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n704_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n506_), .A2(new_n705_), .A3(new_n710_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n666_), .B2(new_n709_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n718_), .A2(KEYINPUT109), .A3(new_n719_), .A4(new_n704_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n457_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n702_), .B1(new_n721_), .B2(new_n213_), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n701_), .A2(new_n214_), .A3(new_n406_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n701_), .A2(new_n214_), .A3(new_n406_), .A4(new_n724_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n714_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n718_), .B2(new_n704_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n719_), .A2(KEYINPUT109), .ZN(new_n731_));
  AOI211_X1 g530(.A(new_n703_), .B(new_n731_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n406_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n728_), .B1(new_n733_), .B2(G36gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n726_), .A2(new_n727_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n497_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n214_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT46), .B1(new_n740_), .B2(KEYINPUT112), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1329gat));
  NAND3_X1  g541(.A1(new_n701_), .A2(new_n212_), .A3(new_n466_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n500_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(new_n212_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1330gat));
  NAND3_X1  g546(.A1(new_n701_), .A2(new_n209_), .A3(new_n352_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n495_), .B1(new_n715_), .B2(new_n720_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n209_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1331gat));
  NOR3_X1   g551(.A1(new_n666_), .A2(new_n590_), .A3(new_n255_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n753_), .A2(new_n605_), .A3(new_n709_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n456_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n668_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(KEYINPUT114), .A3(new_n668_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n456_), .A2(G57gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n760_), .B2(new_n761_), .ZN(G1332gat));
  INV_X1    g561(.A(G64gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n754_), .A2(new_n763_), .A3(new_n406_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n406_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G64gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n766_), .A2(new_n767_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n754_), .A2(new_n771_), .A3(new_n466_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n758_), .A2(new_n466_), .A3(new_n759_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G71gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G71gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT116), .B(new_n772_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1334gat));
  NAND3_X1  g580(.A1(new_n754_), .A2(new_n511_), .A3(new_n352_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n760_), .A2(new_n352_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G78gat), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(KEYINPUT50), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(KEYINPUT50), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(G1335gat));
  NOR4_X1   g586(.A1(new_n700_), .A2(new_n666_), .A3(new_n590_), .A4(new_n255_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n456_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n590_), .A2(new_n255_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n718_), .A2(new_n604_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n456_), .A2(G85gat), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT117), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n789_), .A2(G85gat), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT118), .ZN(G1336gat));
  AOI21_X1  g594(.A(G92gat), .B1(new_n788_), .B2(new_n406_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n791_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n406_), .A2(G92gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(G1337gat));
  NAND3_X1  g598(.A1(new_n788_), .A2(new_n550_), .A3(new_n466_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT119), .ZN(new_n801_));
  INV_X1    g600(.A(G99gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n797_), .B2(new_n466_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n788_), .A2(new_n551_), .A3(new_n352_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n718_), .A2(new_n604_), .A3(new_n352_), .A4(new_n790_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(G106gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n808_), .B2(G106gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n407_), .A2(new_n456_), .A3(new_n466_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n255_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n709_), .A2(new_n605_), .A3(new_n590_), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(KEYINPUT54), .C1(new_n645_), .C2(new_n255_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT55), .B1(new_n569_), .B2(new_n571_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n570_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n548_), .A2(new_n556_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n507_), .B1(new_n566_), .B2(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n824_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n823_), .B1(new_n829_), .B2(new_n581_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n572_), .A2(new_n825_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n826_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n828_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n579_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(KEYINPUT121), .B(new_n823_), .C1(new_n829_), .C2(new_n581_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n255_), .A2(new_n837_), .A3(new_n582_), .A4(new_n838_), .ZN(new_n839_));
  AND4_X1   g638(.A1(new_n242_), .A2(new_n232_), .A3(new_n236_), .A4(new_n238_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n233_), .B2(new_n241_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n253_), .B1(new_n841_), .B2(new_n249_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n583_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n667_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT57), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n830_), .A2(new_n835_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n582_), .A3(new_n842_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n849_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n847_), .A2(new_n582_), .A3(new_n842_), .A4(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n850_), .A2(new_n707_), .A3(new_n708_), .A4(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n844_), .B2(KEYINPUT57), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n604_), .B1(new_n846_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n814_), .B1(new_n822_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n255_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(KEYINPUT123), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n853_), .B(new_n859_), .C1(new_n844_), .C2(KEYINPUT57), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n858_), .A2(new_n845_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n821_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n820_), .B1(new_n816_), .B2(KEYINPUT54), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n861_), .A2(new_n604_), .B1(new_n864_), .B2(new_n819_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(KEYINPUT59), .A3(new_n814_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n856_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n815_), .A2(new_n416_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n857_), .B1(new_n869_), .B2(new_n870_), .ZN(G1340gat));
  OAI21_X1  g670(.A(new_n408_), .B1(new_n590_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n856_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n408_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n866_), .A2(new_n590_), .A3(new_n868_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n408_), .ZN(G1341gat));
  AOI21_X1  g674(.A(G127gat), .B1(new_n856_), .B2(new_n605_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n605_), .A2(G127gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT124), .Z(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n869_), .B2(new_n878_), .ZN(G1342gat));
  AOI21_X1  g678(.A(G134gat), .B1(new_n856_), .B2(new_n667_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n710_), .A2(G134gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n869_), .B2(new_n881_), .ZN(G1343gat));
  AOI21_X1  g681(.A(new_n466_), .B1(new_n822_), .B2(new_n855_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n495_), .A2(new_n406_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n456_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n815_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n257_), .ZN(G1344gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n590_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n258_), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n885_), .A2(new_n604_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  NOR3_X1   g691(.A1(new_n885_), .A2(new_n633_), .A3(new_n709_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n883_), .A2(new_n456_), .A3(new_n667_), .A4(new_n884_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n633_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT125), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n897_), .A3(new_n633_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n893_), .B1(new_n896_), .B2(new_n898_), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n497_), .A2(new_n456_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n901_), .A2(new_n352_), .A3(new_n500_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n861_), .A2(new_n604_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n822_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n246_), .B1(new_n905_), .B2(new_n255_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n361_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n865_), .A2(new_n815_), .A3(new_n907_), .A4(new_n903_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT62), .B1(new_n906_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n865_), .A2(new_n815_), .A3(new_n903_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n246_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1348gat));
  INV_X1    g712(.A(new_n590_), .ZN(new_n914_));
  AOI21_X1  g713(.A(G176gat), .B1(new_n905_), .B2(new_n914_), .ZN(new_n915_));
  AOI211_X1 g714(.A(new_n355_), .B(new_n590_), .C1(new_n822_), .C2(new_n855_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n902_), .B2(new_n916_), .ZN(G1349gat));
  NOR2_X1   g716(.A1(new_n604_), .A2(new_n372_), .ZN(new_n918_));
  INV_X1    g717(.A(G183gat), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n864_), .A2(new_n605_), .A3(new_n819_), .A4(new_n902_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n905_), .A2(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n905_), .A2(new_n667_), .A3(new_n373_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n904_), .A2(new_n822_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n710_), .A3(new_n902_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n924_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT126), .B1(new_n924_), .B2(G190gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n922_), .B1(new_n925_), .B2(new_n926_), .ZN(G1351gat));
  NAND4_X1  g726(.A1(new_n883_), .A2(new_n255_), .A3(new_n352_), .A4(new_n900_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g728(.A1(new_n883_), .A2(new_n900_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n930_), .A2(new_n914_), .A3(new_n352_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G204gat), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n930_), .A2(new_n309_), .A3(new_n914_), .A4(new_n352_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1353gat));
  AOI21_X1  g733(.A(new_n604_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT127), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n883_), .A2(new_n352_), .A3(new_n900_), .A4(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n937_), .B(new_n938_), .Z(G1354gat));
  AND2_X1   g738(.A1(new_n930_), .A2(new_n352_), .ZN(new_n940_));
  INV_X1    g739(.A(G218gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n709_), .A2(new_n941_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n930_), .A2(new_n667_), .A3(new_n352_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n940_), .A2(new_n942_), .B1(new_n943_), .B2(new_n941_), .ZN(G1355gat));
endmodule


