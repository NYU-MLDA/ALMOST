//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n206_));
  AND3_X1   g005(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n211_), .A2(new_n202_), .A3(new_n203_), .A4(new_n204_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G85gat), .B(G92gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n217_), .A3(new_n214_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  AOI211_X1 g024(.A(new_n208_), .B(new_n207_), .C1(new_n225_), .C2(new_n204_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n216_), .A2(new_n218_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT69), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n228_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n235_), .A3(KEYINPUT15), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n235_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT15), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n227_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT34), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n226_), .A2(new_n224_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n218_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n217_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n246_), .B1(new_n250_), .B2(new_n237_), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n240_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G190gat), .B(G218gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G134gat), .B(G162gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(KEYINPUT36), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n245_), .B1(new_n240_), .B2(new_n251_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n252_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n255_), .B(KEYINPUT36), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n258_), .A2(new_n261_), .A3(KEYINPUT37), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT37), .B1(new_n258_), .B2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G127gat), .B(G155gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G183gat), .B(G211gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT70), .ZN(new_n272_));
  INV_X1    g071(.A(G15gat), .ZN(new_n273_));
  INV_X1    g072(.A(G22gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G15gat), .A2(G22gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G1gat), .A2(G8gat), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n275_), .A2(new_n276_), .B1(KEYINPUT14), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n272_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G64gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G57gat), .ZN(new_n283_));
  INV_X1    g082(.A(G57gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G64gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n285_), .A3(KEYINPUT11), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT66), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n285_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT11), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n283_), .A2(new_n285_), .A3(new_n291_), .A4(KEYINPUT11), .ZN(new_n292_));
  AND2_X1   g091(.A1(G71gat), .A2(G78gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G71gat), .A2(G78gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n287_), .A2(new_n290_), .A3(new_n292_), .A4(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n287_), .A2(new_n292_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n281_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n281_), .A2(new_n299_), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT72), .B(KEYINPUT17), .Z(new_n302_));
  OR4_X1    g101(.A1(new_n270_), .A2(new_n300_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n270_), .B(KEYINPUT17), .Z(new_n304_));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G57gat), .B(G64gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n295_), .B1(new_n307_), .B2(KEYINPUT11), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n291_), .B1(new_n307_), .B2(KEYINPUT11), .ZN(new_n309_));
  AND4_X1   g108(.A1(new_n291_), .A2(new_n283_), .A3(new_n285_), .A4(KEYINPUT11), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n296_), .A3(KEYINPUT67), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT73), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n304_), .B1(new_n314_), .B2(new_n281_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n281_), .B2(new_n314_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n303_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n265_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT12), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n311_), .A2(new_n296_), .A3(KEYINPUT67), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT67), .B1(new_n311_), .B2(new_n296_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n323_), .B2(new_n227_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G230gat), .A2(G233gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n216_), .A2(new_n218_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n306_), .A2(new_n326_), .A3(new_n247_), .A4(new_n312_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n320_), .B1(new_n311_), .B2(new_n296_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n250_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n325_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n327_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n323_), .A2(new_n227_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT5), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G176gat), .B(G204gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n335_), .A2(new_n340_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT13), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n319_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT74), .Z(new_n350_));
  INV_X1    g149(.A(KEYINPUT21), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT80), .B(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(G197gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G211gat), .B(G218gat), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n353_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n351_), .B1(G197gat), .B2(G204gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n354_), .A2(new_n355_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n357_), .A2(KEYINPUT21), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369_));
  INV_X1    g168(.A(G141gat), .ZN(new_n370_));
  INV_X1    g169(.A(G148gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT78), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n372_), .B(new_n373_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n375_), .A2(new_n374_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n367_), .B(new_n368_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n367_), .A2(KEYINPUT1), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(G155gat), .A3(G162gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n381_), .A3(new_n368_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n370_), .A2(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n365_), .B(new_n366_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n356_), .A2(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n378_), .B2(new_n385_), .ZN(new_n390_));
  OAI211_X1 g189(.A(G228gat), .B(G233gat), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT82), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n396_), .A3(new_n393_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n393_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n388_), .A2(new_n391_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT81), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n388_), .A2(new_n391_), .A3(new_n401_), .A4(new_n398_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n395_), .A2(new_n397_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G22gat), .B(G50gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n378_), .A2(new_n385_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT28), .B1(new_n406_), .B2(KEYINPUT29), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n406_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n405_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n407_), .A3(new_n404_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n410_), .A2(new_n412_), .A3(KEYINPUT79), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT79), .B1(new_n410_), .B2(new_n412_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n403_), .A2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n410_), .A2(new_n412_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n394_), .A2(KEYINPUT83), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n394_), .A2(KEYINPUT83), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n399_), .B(new_n417_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n420_), .A3(KEYINPUT84), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n426_));
  INV_X1    g225(.A(G169gat), .ZN(new_n427_));
  INV_X1    g226(.A(G176gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT24), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT23), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT24), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n431_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n437_));
  INV_X1    g236(.A(G183gat), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT25), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT26), .B(G190gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT25), .B1(new_n437_), .B2(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n433_), .B1(G183gat), .B2(G190gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n427_), .A2(new_n428_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G169gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n428_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n436_), .A2(new_n442_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n426_), .B1(new_n447_), .B2(new_n389_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n430_), .B1(new_n429_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n449_), .B2(new_n429_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT25), .B(G183gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n440_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n433_), .A3(new_n435_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n443_), .A2(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n365_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n448_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G226gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT19), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G8gat), .B(G36gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n466_), .A2(new_n467_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n463_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n466_), .A2(new_n467_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n389_), .A2(new_n455_), .A3(new_n454_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT86), .ZN(new_n476_));
  INV_X1    g275(.A(new_n460_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT20), .B(new_n477_), .C1(new_n447_), .C2(new_n389_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n461_), .B(new_n474_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n389_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n456_), .A2(new_n365_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n460_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n448_), .A2(new_n477_), .A3(new_n457_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n471_), .A2(KEYINPUT95), .A3(new_n473_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT95), .B1(new_n471_), .B2(new_n473_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n479_), .A2(new_n488_), .A3(KEYINPUT27), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n479_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n474_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n461_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n481_), .A2(KEYINPUT86), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n475_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n478_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n492_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n496_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n478_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n501_), .A2(KEYINPUT89), .A3(new_n461_), .A4(new_n474_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n491_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT27), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n489_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G127gat), .B(G134gat), .Z(new_n507_));
  XOR2_X1   g306(.A(G113gat), .B(G120gat), .Z(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n386_), .B(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n406_), .A2(new_n509_), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n514_), .A2(KEYINPUT90), .ZN(new_n515_));
  INV_X1    g314(.A(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n386_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n406_), .A2(new_n509_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT4), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(KEYINPUT90), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n515_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n512_), .B1(new_n511_), .B2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G1gat), .B(G29gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT91), .B(G85gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT0), .B(G57gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT94), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n522_), .A2(KEYINPUT94), .A3(new_n528_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G227gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n273_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G43gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G71gat), .B(G99gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n447_), .A2(KEYINPUT30), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n447_), .A2(KEYINPUT30), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n536_), .B(new_n541_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n544_), .A2(KEYINPUT77), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n541_), .A2(new_n536_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n542_), .A2(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n536_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n535_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n535_), .A3(new_n549_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n509_), .A3(new_n552_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n545_), .A2(new_n535_), .A3(new_n549_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n516_), .B1(new_n554_), .B2(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NOR4_X1   g355(.A1(new_n425_), .A2(new_n506_), .A3(new_n534_), .A4(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n416_), .A2(new_n420_), .A3(KEYINPUT84), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT84), .B1(new_n416_), .B2(new_n420_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n505_), .B(new_n533_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT96), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n425_), .A2(new_n562_), .A3(new_n533_), .A4(new_n505_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n564_));
  INV_X1    g363(.A(new_n484_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n474_), .A2(KEYINPUT32), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n484_), .A2(KEYINPUT93), .A3(KEYINPUT32), .A4(new_n474_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n474_), .A2(KEYINPUT92), .A3(KEYINPUT32), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n501_), .A2(new_n461_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(new_n568_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n521_), .A2(new_n511_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n512_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n528_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT33), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n527_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n521_), .B2(new_n511_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n491_), .A2(new_n502_), .A3(new_n498_), .A4(new_n579_), .ZN(new_n580_));
  OAI22_X1  g379(.A1(new_n533_), .A2(new_n573_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n558_), .A2(new_n559_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n561_), .A2(new_n563_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n557_), .B1(new_n584_), .B2(new_n556_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n279_), .A2(new_n237_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n279_), .A2(new_n237_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n279_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n239_), .B2(new_n236_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n587_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(new_n586_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n594_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n585_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n350_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n533_), .A2(G1gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n603_), .B(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n258_), .A2(new_n261_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n585_), .A2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n347_), .A2(new_n318_), .A3(new_n599_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n533_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n606_), .A2(KEYINPUT98), .A3(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(G8gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n601_), .A2(new_n618_), .A3(new_n506_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n611_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n506_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n621_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n619_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT40), .B(new_n619_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(new_n556_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n273_), .B1(new_n620_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n601_), .A2(new_n273_), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n633_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n611_), .B2(new_n582_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n601_), .A2(new_n274_), .A3(new_n425_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1327gat));
  NOR3_X1   g440(.A1(new_n347_), .A2(new_n607_), .A3(new_n317_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n600_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n534_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n264_), .B(KEYINPUT100), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n585_), .B2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n264_), .A2(KEYINPUT43), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT101), .B1(new_n585_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651_));
  AOI22_X1  g450(.A1(KEYINPUT96), .A2(new_n560_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n631_), .B1(new_n652_), .B2(new_n563_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n651_), .B(new_n648_), .C1(new_n653_), .C2(new_n557_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n647_), .A2(new_n650_), .A3(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n347_), .A2(new_n317_), .A3(new_n599_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(G29gat), .A3(new_n534_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n645_), .B1(new_n658_), .B2(new_n661_), .ZN(G1328gat));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n506_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G36gat), .B1(new_n663_), .B2(new_n660_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n505_), .A2(G36gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n643_), .A2(KEYINPUT45), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT45), .B1(new_n643_), .B2(new_n666_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n664_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n664_), .B2(new_n675_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(G1329gat));
  INV_X1    g477(.A(G43gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(new_n643_), .B2(new_n556_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT105), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n657_), .A2(G43gat), .A3(new_n631_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n660_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n681_), .B(new_n685_), .C1(new_n660_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n644_), .B2(new_n425_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n657_), .A2(G50gat), .A3(new_n425_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n661_), .ZN(G1331gat));
  NOR3_X1   g489(.A1(new_n348_), .A2(new_n318_), .A3(new_n598_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n609_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n533_), .A2(new_n284_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT107), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n319_), .A2(new_n347_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n599_), .B1(new_n653_), .B2(new_n557_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT106), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT106), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n534_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n696_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(G1332gat));
  OAI21_X1  g504(.A(G64gat), .B1(new_n692_), .B2(new_n505_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n701_), .A2(new_n282_), .A3(new_n506_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  OAI21_X1  g509(.A(G71gat), .B1(new_n692_), .B2(new_n556_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT49), .ZN(new_n712_));
  INV_X1    g511(.A(new_n701_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n556_), .A2(G71gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1334gat));
  OAI21_X1  g514(.A(G78gat), .B1(new_n692_), .B2(new_n582_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT50), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n582_), .A2(G78gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT110), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n713_), .B2(new_n719_), .ZN(G1335gat));
  NAND3_X1  g519(.A1(new_n347_), .A2(new_n608_), .A3(new_n318_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n221_), .A3(new_n534_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n347_), .A2(new_n318_), .A3(new_n599_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT111), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n655_), .A2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n533_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1336gat));
  AOI21_X1  g527(.A(G92gat), .B1(new_n722_), .B2(new_n506_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n726_), .A2(new_n505_), .A3(new_n220_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1337gat));
  AND2_X1   g530(.A1(new_n631_), .A2(new_n225_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n722_), .A2(new_n732_), .B1(new_n733_), .B2(KEYINPUT51), .ZN(new_n734_));
  OAI21_X1  g533(.A(G99gat), .B1(new_n726_), .B2(new_n556_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n733_), .A2(KEYINPUT51), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n736_), .B(new_n737_), .Z(G1338gat));
  NAND3_X1  g537(.A1(new_n722_), .A2(new_n204_), .A3(new_n425_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n655_), .A2(new_n425_), .A3(new_n725_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G106gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n608_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n592_), .B2(new_n587_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n239_), .A2(new_n236_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT116), .B(new_n588_), .C1(new_n750_), .C2(new_n591_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n749_), .A2(new_n751_), .A3(G229gat), .A4(G233gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n588_), .A2(new_n589_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n597_), .B1(new_n753_), .B2(new_n586_), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n752_), .A2(new_n754_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n755_), .B(new_n758_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n598_), .A2(new_n341_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n330_), .A2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n327_), .A2(new_n329_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(KEYINPUT55), .A3(new_n325_), .A4(new_n324_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n327_), .A2(new_n329_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT12), .B1(new_n313_), .B2(new_n250_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n331_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(new_n765_), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT113), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n769_), .A2(new_n339_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n771_), .B1(new_n769_), .B2(new_n339_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n339_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n773_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n761_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n760_), .B1(new_n780_), .B2(KEYINPUT115), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n769_), .A2(new_n339_), .A3(new_n774_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n769_), .A2(new_n339_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n772_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n598_), .A2(new_n341_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT115), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n747_), .B1(new_n781_), .B2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n755_), .A2(new_n341_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n339_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n778_), .A2(KEYINPUT118), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n790_), .B(new_n793_), .C1(new_n794_), .C2(new_n791_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT58), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n264_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n789_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n785_), .A2(new_n786_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n787_), .A3(new_n760_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n607_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n318_), .B1(new_n801_), .B2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n319_), .A2(new_n599_), .A3(new_n348_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT54), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n425_), .A2(new_n506_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n534_), .A3(new_n631_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT120), .B1(new_n801_), .B2(new_n806_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n607_), .B1(new_n781_), .B2(new_n788_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n746_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n805_), .A2(new_n747_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n318_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n813_), .B1(new_n822_), .B2(new_n809_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n815_), .B1(new_n823_), .B2(new_n811_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT121), .B(new_n815_), .C1(new_n823_), .C2(new_n811_), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n599_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n823_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n831_), .B2(new_n599_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1340gat));
  OAI21_X1  g632(.A(G120gat), .B1(new_n824_), .B2(new_n348_), .ZN(new_n834_));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n348_), .B2(KEYINPUT60), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(KEYINPUT60), .B2(new_n835_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n834_), .B1(new_n831_), .B2(new_n837_), .ZN(G1341gat));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n318_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n826_), .A2(new_n827_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n831_), .B2(new_n318_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n264_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n826_), .A2(new_n827_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n831_), .B2(new_n607_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1343gat));
  NAND2_X1  g647(.A1(new_n822_), .A2(new_n809_), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n631_), .A2(new_n582_), .A3(new_n506_), .A4(new_n533_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n599_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT122), .B(G141gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n851_), .A2(new_n348_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n371_), .ZN(G1345gat));
  NOR2_X1   g655(.A1(new_n851_), .A2(new_n318_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT61), .B(G155gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n851_), .B2(new_n607_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n851_), .A2(new_n860_), .A3(new_n646_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT123), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n861_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1347gat));
  NOR4_X1   g667(.A1(new_n425_), .A2(new_n534_), .A3(new_n556_), .A4(new_n505_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n810_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870_), .B2(new_n599_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(KEYINPUT62), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(KEYINPUT62), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n598_), .A2(new_n445_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(KEYINPUT124), .Z(new_n875_));
  OAI22_X1  g674(.A1(new_n872_), .A2(new_n873_), .B1(new_n870_), .B2(new_n875_), .ZN(G1348gat));
  NAND2_X1  g675(.A1(new_n849_), .A2(new_n869_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n348_), .A2(new_n428_), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n878_), .A2(KEYINPUT125), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT125), .B1(new_n878_), .B2(new_n879_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n870_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G176gat), .B1(new_n882_), .B2(new_n347_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n880_), .A2(new_n881_), .A3(new_n883_), .ZN(G1349gat));
  OAI21_X1  g683(.A(new_n438_), .B1(new_n877_), .B2(new_n318_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n318_), .A2(new_n452_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n810_), .A2(new_n869_), .A3(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT126), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT127), .B1(new_n886_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n889_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT127), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n885_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n870_), .B2(new_n264_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n608_), .A2(new_n440_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n870_), .B2(new_n896_), .ZN(G1351gat));
  NAND2_X1  g696(.A1(new_n425_), .A2(new_n533_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n506_), .A2(new_n556_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n898_), .B(new_n899_), .C1(new_n822_), .C2(new_n809_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n598_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n347_), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n352_), .B(G204gat), .S(new_n903_), .Z(G1353gat));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n317_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  INV_X1    g708(.A(G218gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n900_), .A2(new_n910_), .A3(new_n608_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n900_), .A2(new_n265_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n910_), .ZN(G1355gat));
endmodule


