//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204_));
  OAI22_X1  g003(.A1(new_n204_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .A4(KEYINPUT86), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  OAI22_X1  g009(.A1(new_n207_), .A2(new_n208_), .B1(new_n210_), .B2(KEYINPUT87), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(KEYINPUT87), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n205_), .B(new_n209_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT88), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n202_), .B(new_n203_), .C1(new_n213_), .C2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G155gat), .A3(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT85), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n203_), .A4(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n222_), .C1(new_n220_), .C2(new_n219_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT28), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n224_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G22gat), .B(G50gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n227_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n231_), .B2(new_n225_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT92), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n235_));
  XOR2_X1   g034(.A(G211gat), .B(G218gat), .Z(new_n236_));
  OAI22_X1  g035(.A1(new_n235_), .A2(new_n236_), .B1(KEYINPUT21), .B2(new_n234_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n239_), .B1(KEYINPUT29), .B2(new_n224_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT89), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n239_), .B2(KEYINPUT91), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n240_), .A2(new_n243_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n229_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n231_), .A2(new_n225_), .A3(new_n228_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n233_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n252_));
  OAI221_X1 g051(.A(KEYINPUT92), .B1(new_n230_), .B2(new_n232_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G78gat), .B(G106gat), .Z(new_n254_));
  AND3_X1   g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT27), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  INV_X1    g059(.A(G183gat), .ZN(new_n261_));
  INV_X1    g060(.A(G190gat), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT23), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT23), .B1(new_n261_), .B2(new_n262_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT79), .B(G190gat), .Z(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(G183gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT83), .B(G176gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT22), .B(G169gat), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n269_), .A2(new_n270_), .B1(G169gat), .B2(G176gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT82), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n265_), .B(KEYINPUT81), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n264_), .ZN(new_n276_));
  OR2_X1    g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT24), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT25), .B(G183gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT80), .B(KEYINPUT26), .Z(new_n283_));
  OAI221_X1 g082(.A(new_n281_), .B1(new_n267_), .B2(new_n282_), .C1(new_n262_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n277_), .A2(KEYINPUT24), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n280_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n276_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n273_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n260_), .B1(new_n290_), .B2(new_n239_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n239_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT26), .B(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n281_), .A2(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n297_), .A2(KEYINPUT93), .A3(new_n286_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT93), .B1(new_n297_), .B2(new_n286_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n266_), .B(new_n279_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n265_), .A2(KEYINPUT81), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n265_), .A2(KEYINPUT81), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n263_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n271_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT94), .B1(new_n295_), .B2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n295_), .A2(KEYINPUT94), .A3(new_n306_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n291_), .B(new_n294_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT20), .B1(new_n295_), .B2(new_n306_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT95), .B1(new_n290_), .B2(new_n239_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT82), .B1(new_n303_), .B2(new_n278_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n289_), .A2(new_n312_), .A3(new_n286_), .A4(new_n284_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n272_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n295_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n310_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n309_), .B1(new_n317_), .B2(new_n294_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G64gat), .B(G92gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT97), .ZN(new_n320_));
  XOR2_X1   g119(.A(G8gat), .B(G36gat), .Z(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n259_), .B1(new_n318_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT102), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n308_), .A2(new_n307_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n295_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n293_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n310_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n315_), .B1(new_n314_), .B2(new_n295_), .ZN(new_n332_));
  AOI211_X1 g131(.A(KEYINPUT95), .B(new_n239_), .C1(new_n313_), .C2(new_n272_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n294_), .B(new_n331_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n327_), .B1(new_n335_), .B2(new_n325_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(new_n334_), .A3(KEYINPUT102), .A4(new_n324_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n326_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341_));
  XOR2_X1   g140(.A(G113gat), .B(G120gat), .Z(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND3_X1  g142(.A1(new_n224_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT99), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT99), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n339_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n216_), .A2(KEYINPUT98), .A3(new_n223_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n349_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT4), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT100), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n347_), .A2(KEYINPUT100), .A3(new_n353_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n352_), .A2(new_n339_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n356_), .A2(new_n361_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n354_), .A2(new_n355_), .B1(new_n352_), .B2(new_n339_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n361_), .B1(new_n366_), .B2(new_n362_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n335_), .A2(new_n325_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n324_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n259_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n258_), .A2(new_n338_), .A3(new_n368_), .A4(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(new_n370_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n339_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n345_), .A2(new_n346_), .B1(G225gat), .B2(G233gat), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n361_), .B(new_n374_), .C1(new_n375_), .C2(new_n353_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n364_), .B2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n366_), .A2(KEYINPUT33), .A3(new_n361_), .A4(new_n362_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n335_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n318_), .A2(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n382_), .B(new_n383_), .C1(new_n365_), .C2(new_n367_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n372_), .B1(new_n385_), .B2(new_n258_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT84), .B(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n314_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(new_n343_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(G15gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT30), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT31), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n338_), .A2(new_n257_), .A3(new_n371_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT103), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n338_), .A2(new_n257_), .A3(KEYINPUT103), .A4(new_n371_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n368_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n386_), .A2(new_n400_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G1gat), .A2(G8gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT14), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT73), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n413_), .A3(KEYINPUT14), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G15gat), .B(G22gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G1gat), .B(G8gat), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n417_), .A2(new_n412_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G43gat), .B(G50gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G36gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G29gat), .ZN(new_n425_));
  INV_X1    g224(.A(G29gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G36gat), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(new_n427_), .A3(KEYINPUT68), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT68), .B1(new_n425_), .B2(new_n427_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n423_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n427_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n425_), .A2(new_n427_), .A3(KEYINPUT68), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n422_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n421_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n421_), .A2(new_n436_), .A3(KEYINPUT76), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n430_), .A2(new_n435_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(KEYINPUT75), .A3(new_n419_), .A4(new_n420_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT75), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n421_), .B2(new_n436_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT77), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT77), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n441_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT15), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n436_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n421_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n446_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n449_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n453_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n409_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n453_), .A2(new_n458_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n461_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT78), .A3(new_n463_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G190gat), .B(G218gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G134gat), .B(G162gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n474_), .B(KEYINPUT36), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n477_));
  AND3_X1   g276(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT9), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G85gat), .B(G92gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n481_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT10), .B(G99gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(G106gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT64), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n492_), .A2(new_n493_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT64), .ZN(new_n495_));
  NOR2_X1   g294(.A1(G85gat), .A2(G92gat), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n485_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT9), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n494_), .A2(new_n495_), .A3(new_n480_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n489_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n501_));
  INV_X1    g300(.A(G99gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n493_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n503_), .A2(new_n506_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n485_), .A2(new_n496_), .A3(KEYINPUT8), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(KEYINPUT65), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  INV_X1    g315(.A(new_n508_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT66), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n503_), .A2(new_n520_), .A3(new_n508_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n480_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n516_), .B1(new_n522_), .B2(new_n497_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n500_), .B(new_n442_), .C1(new_n515_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n506_), .A2(new_n507_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n503_), .A2(new_n508_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(KEYINPUT66), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n482_), .B1(new_n529_), .B2(new_n521_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n513_), .B(new_n514_), .C1(new_n530_), .C2(new_n516_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n531_), .A2(KEYINPUT69), .A3(new_n442_), .A4(new_n500_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT34), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n500_), .B1(new_n515_), .B2(new_n523_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n455_), .A2(new_n540_), .B1(new_n537_), .B2(new_n536_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n533_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n533_), .B2(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n477_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n538_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n533_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(KEYINPUT71), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n476_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT70), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n542_), .A2(new_n543_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n474_), .A2(KEYINPUT36), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  AND4_X1   g352(.A1(new_n550_), .A2(new_n546_), .A3(new_n552_), .A4(new_n547_), .ZN(new_n554_));
  OAI22_X1  g353(.A1(new_n549_), .A2(KEYINPUT72), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556_));
  AOI211_X1 g355(.A(new_n556_), .B(new_n476_), .C1(new_n544_), .C2(new_n548_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n471_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n500_), .B(new_n566_), .C1(new_n515_), .C2(new_n523_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  INV_X1    g369(.A(new_n566_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n540_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n540_), .B2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n568_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n522_), .A2(new_n497_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT8), .ZN(new_n577_));
  INV_X1    g376(.A(new_n514_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT65), .B1(new_n509_), .B2(new_n510_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n577_), .A2(new_n580_), .B1(new_n489_), .B2(new_n499_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n566_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n567_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n575_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n574_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n574_), .B2(new_n584_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n559_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT67), .A3(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n595_), .A3(KEYINPUT13), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT37), .B1(new_n551_), .B2(new_n476_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n551_), .A2(new_n552_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT70), .ZN(new_n603_));
  INV_X1    g402(.A(new_n554_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n601_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n421_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n571_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n610_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  MUX2_X1   g415(.A(new_n615_), .B(KEYINPUT17), .S(new_n614_), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n558_), .A2(new_n600_), .A3(new_n606_), .A4(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n408_), .A2(new_n470_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(G1gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n406_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT38), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n542_), .A2(new_n543_), .A3(new_n477_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT71), .B1(new_n546_), .B2(new_n547_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n475_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n556_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n603_), .A2(new_n604_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n549_), .A2(KEYINPUT72), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n408_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n470_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n600_), .A4(new_n620_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n368_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n624_), .A2(new_n625_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n626_), .A2(new_n638_), .A3(new_n639_), .ZN(G1324gat));
  NAND2_X1  g439(.A1(new_n338_), .A2(new_n371_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G8gat), .B1(new_n637_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT39), .ZN(new_n644_));
  INV_X1    g443(.A(G8gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n622_), .A2(new_n645_), .A3(new_n641_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n637_), .B2(new_n400_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT41), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n622_), .A2(new_n393_), .A3(new_n399_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1326gat));
  OAI21_X1  g451(.A(G22gat), .B1(new_n637_), .B2(new_n257_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n622_), .A2(new_n655_), .A3(new_n258_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n408_), .A2(new_n470_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n600_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(new_n620_), .A3(new_n633_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n406_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n605_), .B1(new_n633_), .B2(new_n471_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n405_), .A2(new_n407_), .ZN(new_n666_));
  AND4_X1   g465(.A1(new_n258_), .A2(new_n338_), .A3(new_n368_), .A4(new_n371_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n258_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n400_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n664_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n408_), .C2(new_n665_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n671_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n659_), .A2(new_n470_), .A3(new_n620_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n426_), .B(new_n368_), .C1(new_n677_), .C2(KEYINPUT44), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n663_), .B1(new_n678_), .B2(new_n680_), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n662_), .A2(new_n424_), .A3(new_n641_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n682_), .B(new_n683_), .Z(new_n684_));
  AOI21_X1  g483(.A(new_n642_), .B1(new_n677_), .B2(KEYINPUT44), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n680_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT46), .B(new_n684_), .C1(new_n686_), .C2(new_n424_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n424_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n684_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n691_), .ZN(G1329gat));
  XOR2_X1   g491(.A(KEYINPUT106), .B(G43gat), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n661_), .B2(new_n400_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n677_), .A2(KEYINPUT44), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(G43gat), .A3(new_n399_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(new_n679_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g497(.A1(new_n661_), .A2(G50gat), .A3(new_n257_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n695_), .A2(new_n258_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n679_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G50gat), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n701_), .A2(new_n700_), .A3(new_n679_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n600_), .A2(new_n636_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n408_), .A2(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n558_), .A2(new_n620_), .A3(new_n606_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n406_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n635_), .A2(new_n620_), .A3(new_n706_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n368_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1332gat));
  OAI21_X1  g514(.A(G64gat), .B1(new_n713_), .B2(new_n642_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT48), .ZN(new_n717_));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n710_), .A2(new_n718_), .A3(new_n641_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n713_), .B2(new_n400_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT49), .ZN(new_n722_));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n710_), .A2(new_n723_), .A3(new_n399_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n713_), .B2(new_n257_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n257_), .A2(G78gat), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT109), .Z(new_n730_));
  NAND2_X1  g529(.A1(new_n710_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n633_), .A2(new_n620_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n708_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G85gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n406_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n707_), .A2(new_n620_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n675_), .A2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(new_n406_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n740_), .B2(new_n736_), .ZN(G1336gat));
  INV_X1    g540(.A(G92gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n734_), .B2(new_n642_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT110), .Z(new_n744_));
  NOR2_X1   g543(.A1(new_n642_), .A2(new_n742_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n739_), .B2(new_n745_), .ZN(G1337gat));
  AOI21_X1  g545(.A(new_n502_), .B1(new_n739_), .B2(new_n399_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n734_), .A2(new_n400_), .A3(new_n487_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n747_), .A2(KEYINPUT111), .A3(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g549(.A1(new_n735_), .A2(new_n493_), .A3(new_n258_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n675_), .A2(new_n258_), .A3(new_n738_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n675_), .A2(KEYINPUT112), .A3(new_n258_), .A4(new_n738_), .ZN(new_n756_));
  AND4_X1   g555(.A1(new_n752_), .A2(new_n755_), .A3(G106gat), .A4(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n493_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n752_), .B1(new_n758_), .B2(new_n756_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n751_), .C1(new_n757_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT59), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n709_), .A2(new_n767_), .A3(new_n470_), .A4(new_n600_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT54), .B1(new_n621_), .B2(new_n636_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT55), .B(new_n569_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n567_), .A2(new_n568_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT12), .B1(new_n581_), .B2(new_n566_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n540_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n774_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n568_), .B1(new_n778_), .B2(new_n567_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT56), .B(new_n588_), .C1(new_n777_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n567_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n575_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n776_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n574_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n785_), .A3(new_n771_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n588_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n781_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n450_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n462_), .B1(new_n457_), .B2(new_n449_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n791_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n452_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n451_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n449_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n796_), .A3(KEYINPUT116), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n468_), .A2(new_n792_), .A3(new_n797_), .A4(new_n590_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n770_), .B1(new_n788_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n588_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n780_), .ZN(new_n803_));
  AND4_X1   g602(.A1(new_n468_), .A2(new_n797_), .A3(new_n792_), .A4(new_n590_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n799_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT117), .B1(new_n665_), .B2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n803_), .A2(KEYINPUT58), .A3(new_n804_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT58), .B1(new_n803_), .B2(new_n804_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n558_), .A2(new_n606_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n468_), .A2(new_n797_), .A3(new_n792_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n596_), .A2(new_n815_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT114), .B(KEYINPUT56), .Z(new_n817_));
  NAND2_X1  g616(.A1(new_n800_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n800_), .A2(KEYINPUT115), .A3(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n780_), .A3(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n466_), .A2(new_n469_), .A3(new_n590_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n814_), .B1(new_n824_), .B2(new_n634_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n466_), .A2(new_n469_), .A3(new_n590_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n821_), .A2(new_n780_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n820_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n633_), .C1(new_n828_), .C2(new_n816_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n807_), .A2(new_n813_), .A3(new_n825_), .A4(new_n829_), .ZN(new_n830_));
  AOI221_X4 g629(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .C1(new_n830_), .C2(new_n619_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n807_), .A2(new_n813_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n825_), .A2(new_n829_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n619_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n768_), .A2(new_n769_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT118), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n831_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n400_), .A2(new_n368_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n405_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n765_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n665_), .A2(new_n806_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n619_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n835_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(KEYINPUT119), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n844_), .B2(new_n845_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT120), .B1(new_n841_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n848_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n846_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n831_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n852_), .B(new_n853_), .C1(new_n854_), .C2(new_n765_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n636_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G113gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n854_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n470_), .A2(G113gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(G1340gat));
  NOR2_X1   g659(.A1(new_n600_), .A2(KEYINPUT60), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  MUX2_X1   g661(.A(KEYINPUT60), .B(new_n861_), .S(new_n862_), .Z(new_n863_));
  NAND2_X1  g662(.A1(new_n854_), .A2(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n841_), .A2(new_n849_), .A3(new_n600_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n862_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT121), .B(new_n864_), .C1(new_n865_), .C2(new_n862_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n619_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n850_), .A2(new_n855_), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n858_), .B2(new_n619_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n873_), .A2(KEYINPUT122), .A3(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1342gat));
  NAND3_X1  g678(.A1(new_n850_), .A2(new_n811_), .A3(new_n855_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G134gat), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n633_), .A2(G134gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n858_), .B2(new_n882_), .ZN(G1343gat));
  NAND2_X1  g682(.A1(new_n834_), .A2(new_n835_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n766_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n834_), .A2(KEYINPUT118), .A3(new_n835_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n399_), .A3(new_n257_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(new_n406_), .A3(new_n642_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n470_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n207_), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n600_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n208_), .ZN(G1345gat));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n619_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT61), .B(G155gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n889_), .A2(new_n897_), .A3(new_n665_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n889_), .B2(new_n633_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT123), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n901_), .B(new_n897_), .C1(new_n889_), .C2(new_n633_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n898_), .B1(new_n900_), .B2(new_n902_), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n642_), .A2(new_n406_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n844_), .A2(new_n399_), .A3(new_n257_), .A4(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n470_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OAI21_X1  g706(.A(G169gat), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n907_), .B2(new_n906_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n910_));
  OR2_X1    g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(new_n270_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n910_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(G1348gat));
  OAI21_X1  g713(.A(new_n269_), .B1(new_n905_), .B2(new_n600_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT126), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n887_), .A2(new_n258_), .ZN(new_n917_));
  AND4_X1   g716(.A1(G176gat), .A2(new_n904_), .A3(new_n399_), .A4(new_n659_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1349gat));
  NOR3_X1   g718(.A1(new_n905_), .A2(new_n281_), .A3(new_n619_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n917_), .A2(new_n399_), .A3(new_n620_), .A4(new_n904_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n261_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n905_), .B2(new_n665_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT127), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n634_), .A2(new_n296_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n905_), .B2(new_n925_), .ZN(G1351gat));
  NAND2_X1  g725(.A1(new_n888_), .A2(new_n904_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n470_), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n600_), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n930_), .B(G204gat), .Z(G1353gat));
  OR2_X1    g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT63), .B(G211gat), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n927_), .A2(new_n619_), .ZN(new_n934_));
  MUX2_X1   g733(.A(new_n932_), .B(new_n933_), .S(new_n934_), .Z(G1354gat));
  OAI21_X1  g734(.A(G218gat), .B1(new_n927_), .B2(new_n665_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n633_), .A2(G218gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n927_), .B2(new_n937_), .ZN(G1355gat));
endmodule


