//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_;
  INV_X1    g000(.A(G127gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G127gat), .A2(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G113gat), .ZN(new_n208_));
  INV_X1    g007(.A(G113gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G120gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n208_), .A2(new_n210_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT87), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(new_n206_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n213_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT31), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G71gat), .B(G99gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT84), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G227gat), .A2(G233gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT85), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n222_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G15gat), .B(G43gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n225_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT26), .B(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT83), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT23), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n238_), .A2(KEYINPUT24), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n235_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT30), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G169gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n237_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n247_), .A3(new_n240_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n244_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n229_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n248_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT30), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(KEYINPUT86), .A3(new_n249_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n228_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT86), .B1(new_n254_), .B2(new_n249_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n225_), .B(new_n226_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n220_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n250_), .A2(new_n251_), .A3(new_n229_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n261_), .B2(new_n257_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n220_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n252_), .A2(new_n228_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n260_), .A2(new_n265_), .A3(KEYINPUT88), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT88), .B1(new_n260_), .B2(new_n265_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G228gat), .A2(G233gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT90), .Z(new_n270_));
  AND2_X1   g069(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(G204gat), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  INV_X1    g073(.A(G204gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G197gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n275_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(G197gat), .B2(G204gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT92), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT92), .B1(new_n279_), .B2(new_n280_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n277_), .B(new_n278_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n276_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n278_), .A2(new_n274_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT93), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(KEYINPUT93), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294_));
  INV_X1    g093(.A(G141gat), .ZN(new_n295_));
  INV_X1    g094(.A(G148gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G155gat), .ZN(new_n304_));
  INV_X1    g103(.A(G162gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(KEYINPUT89), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT89), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(G155gat), .B2(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n303_), .A2(new_n306_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT1), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n311_), .A2(new_n306_), .A3(new_n308_), .A4(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n295_), .A2(new_n296_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n298_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT29), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n270_), .B1(new_n293_), .B2(new_n319_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n317_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT28), .B1(new_n317_), .B2(KEYINPUT29), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G22gat), .B(G50gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n323_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n288_), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n328_), .A2(new_n270_), .A3(new_n319_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n320_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n327_), .B1(new_n320_), .B2(new_n329_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n268_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n290_), .A2(new_n248_), .A3(new_n243_), .A4(new_n291_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n248_), .A2(KEYINPUT94), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n245_), .A2(new_n338_), .A3(new_n247_), .A4(new_n240_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n242_), .A2(new_n232_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n341_), .B2(new_n288_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT19), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n335_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n340_), .A2(new_n248_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n336_), .B1(new_n328_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n292_), .B2(new_n253_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n284_), .A2(KEYINPUT93), .A3(new_n287_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT93), .B1(new_n284_), .B2(new_n287_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n349_), .B(new_n253_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n348_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n346_), .B1(new_n355_), .B2(new_n344_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G64gat), .B(G92gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT101), .B1(new_n356_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT101), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n253_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT95), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n353_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n345_), .B1(new_n368_), .B2(new_n348_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n364_), .B(new_n365_), .C1(new_n369_), .C2(new_n346_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT20), .B(new_n345_), .C1(new_n341_), .C2(new_n288_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n367_), .B2(new_n353_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n345_), .B1(new_n335_), .B2(new_n342_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n362_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n363_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT99), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n219_), .A2(new_n377_), .A3(new_n378_), .A4(new_n317_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n317_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(new_n377_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n317_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n217_), .A2(new_n213_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n382_), .A2(KEYINPUT98), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT98), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n219_), .A2(new_n387_), .A3(new_n317_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n379_), .B(new_n381_), .C1(new_n389_), .C2(new_n378_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n380_), .A3(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393_));
  INV_X1    g192(.A(G85gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT0), .B(G57gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  NAND2_X1  g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n390_), .A2(new_n399_), .A3(new_n391_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(KEYINPUT102), .A3(new_n400_), .ZN(new_n401_));
  AOI211_X1 g200(.A(KEYINPUT102), .B(new_n399_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n376_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n390_), .A2(KEYINPUT33), .A3(new_n399_), .A4(new_n391_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n379_), .B(new_n380_), .C1(new_n389_), .C2(new_n378_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT100), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n386_), .A2(new_n381_), .A3(new_n388_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n397_), .A3(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n409_), .A2(new_n410_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n406_), .B(new_n408_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n374_), .A2(KEYINPUT97), .A3(new_n361_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n373_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n350_), .A2(new_n354_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n361_), .B(new_n417_), .C1(new_n418_), .C2(new_n371_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n361_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT97), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n415_), .B1(new_n416_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n334_), .B1(new_n405_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n426_), .A3(new_n416_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n419_), .B(KEYINPUT27), .C1(new_n356_), .C2(new_n361_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n333_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n333_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n260_), .A2(new_n265_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT103), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n400_), .A2(KEYINPUT102), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n399_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n436_), .B1(new_n439_), .B2(new_n402_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n401_), .A2(new_n403_), .A3(KEYINPUT103), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n429_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n425_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G113gat), .B(G141gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G169gat), .B(G197gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G229gat), .A2(G233gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(G1gat), .B(G8gat), .Z(new_n449_));
  NAND2_X1  g248(.A1(G1gat), .A2(G8gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT14), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G15gat), .A2(G22gat), .ZN(new_n452_));
  AND2_X1   g251(.A1(G15gat), .A2(G22gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT77), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n451_), .B(new_n456_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n449_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G43gat), .B(G50gat), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT73), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G43gat), .B(G50gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT73), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n464_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n462_), .A2(new_n463_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n455_), .A2(new_n449_), .A3(new_n457_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n459_), .A2(new_n466_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n468_), .A2(new_n469_), .A3(new_n467_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n465_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n473_), .A2(new_n458_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT80), .B1(new_n472_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n472_), .A2(new_n476_), .A3(KEYINPUT80), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n448_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n473_), .A2(new_n458_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n470_), .A2(KEYINPUT15), .A3(new_n466_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n481_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n448_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n472_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n447_), .B1(new_n480_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n479_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(new_n490_), .B2(new_n477_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n485_), .A2(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n448_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n447_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n495_), .A2(KEYINPUT81), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n495_), .B2(KEYINPUT81), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n489_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(KEYINPUT81), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT82), .ZN(new_n501_));
  INV_X1    g300(.A(new_n489_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n495_), .A2(KEYINPUT81), .A3(new_n496_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n444_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G92gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n394_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT64), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT9), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n508_), .A2(KEYINPUT64), .A3(new_n512_), .A4(new_n509_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n508_), .A3(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT65), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  NAND3_X1  g320(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(G99gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT10), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT10), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(G99gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n517_), .A2(new_n523_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n514_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT7), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n533_), .B(KEYINPUT66), .C1(G99gat), .C2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n525_), .B(new_n524_), .C1(new_n535_), .C2(KEYINPUT7), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT65), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n521_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT67), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n535_), .A2(KEYINPUT7), .ZN(new_n544_));
  NOR2_X1   g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n517_), .A2(new_n523_), .B1(new_n546_), .B2(new_n534_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT67), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n508_), .A2(new_n509_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT8), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n520_), .A2(new_n522_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n534_), .B2(new_n546_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT8), .B1(new_n554_), .B2(new_n550_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n532_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n474_), .A2(new_n475_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT75), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n484_), .A2(new_n482_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n514_), .A2(new_n560_), .A3(new_n530_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n514_), .B2(new_n530_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT8), .ZN(new_n564_));
  INV_X1    g363(.A(new_n553_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n538_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n550_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n551_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n541_), .B2(KEYINPUT67), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n570_), .B2(new_n549_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n559_), .B1(new_n563_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n558_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT35), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT75), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n551_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n517_), .A2(new_n523_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n578_), .A2(new_n548_), .A3(new_n538_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n555_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n557_), .A3(new_n531_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT34), .ZN(new_n583_));
  INV_X1    g382(.A(G232gat), .ZN(new_n584_));
  INV_X1    g383(.A(G233gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n558_), .A2(new_n575_), .A3(new_n588_), .A4(new_n572_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n583_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n587_), .B1(new_n583_), .B2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n574_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n586_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(KEYINPUT35), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(KEYINPUT36), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n592_), .A2(new_n596_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT76), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n592_), .A2(new_n596_), .A3(KEYINPUT76), .A4(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n592_), .A2(new_n596_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n599_), .B(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT37), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n612_), .A3(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G57gat), .B(G64gat), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT11), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT11), .ZN(new_n618_));
  XOR2_X1   g417(.A(G71gat), .B(G78gat), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n481_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G127gat), .B(G155gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT16), .B(G183gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT17), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n629_), .B(KEYINPUT17), .Z(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n625_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT78), .Z(new_n634_));
  NOR2_X1   g433(.A1(new_n615_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n622_), .B1(new_n580_), .B2(new_n531_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n531_), .A2(KEYINPUT68), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n514_), .A2(new_n560_), .A3(new_n530_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n555_), .A2(new_n552_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT12), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n622_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n636_), .A2(KEYINPUT12), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT69), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n580_), .A2(new_n531_), .A3(new_n622_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n643_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n622_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n571_), .B2(new_n532_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n646_), .B1(new_n652_), .B2(new_n645_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(new_n275_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT5), .B(G176gat), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n655_), .B(new_n656_), .Z(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n650_), .A2(new_n653_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT70), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT71), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n664_), .B2(KEYINPUT13), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n662_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT72), .Z(new_n669_));
  NAND2_X1  g468(.A1(new_n635_), .A2(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n670_), .A2(KEYINPUT79), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(KEYINPUT79), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n506_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n442_), .A2(G1gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n634_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n444_), .A2(new_n610_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n442_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n668_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n505_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n679_), .A3(new_n682_), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n676_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT38), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n675_), .A2(KEYINPUT104), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT104), .B1(new_n675_), .B2(new_n685_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(G1324gat));
  NAND2_X1  g487(.A1(new_n678_), .A2(new_n682_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G8gat), .B1(new_n689_), .B2(new_n429_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT39), .ZN(new_n691_));
  INV_X1    g490(.A(new_n673_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n429_), .A2(G8gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n694_), .B(new_n696_), .ZN(G1325gat));
  INV_X1    g496(.A(new_n268_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G15gat), .B1(new_n689_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT41), .Z(new_n700_));
  OR2_X1    g499(.A1(new_n698_), .A2(G15gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n692_), .B2(new_n701_), .ZN(G1326gat));
  OAI21_X1  g501(.A(G22gat), .B1(new_n689_), .B2(new_n431_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n431_), .A2(G22gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n692_), .B2(new_n706_), .ZN(G1327gat));
  NAND3_X1  g506(.A1(new_n668_), .A2(new_n634_), .A3(new_n505_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n668_), .A2(KEYINPUT107), .A3(new_n634_), .A4(new_n505_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n611_), .A2(new_n444_), .A3(new_n613_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT43), .B1(new_n713_), .B2(KEYINPUT108), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n712_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(G29gat), .A3(new_n679_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n712_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n610_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n444_), .A2(new_n722_), .A3(new_n634_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n682_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n442_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n719_), .A2(new_n721_), .B1(G29gat), .B2(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT109), .Z(G1328gat));
  AND2_X1   g527(.A1(new_n429_), .A2(KEYINPUT111), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n429_), .A2(KEYINPUT111), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n725_), .A2(G36gat), .A3(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT45), .Z(new_n734_));
  INV_X1    g533(.A(G36gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n429_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT110), .B(new_n735_), .C1(new_n736_), .C2(new_n720_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738_));
  INV_X1    g537(.A(new_n429_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n718_), .A2(new_n739_), .A3(new_n720_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n740_), .B2(G36gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n734_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n734_), .B(KEYINPUT46), .C1(new_n737_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  NAND3_X1  g545(.A1(new_n718_), .A2(G43gat), .A3(new_n433_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n725_), .A2(new_n698_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n747_), .A2(new_n721_), .B1(G43gat), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g549(.A1(new_n718_), .A2(G50gat), .A3(new_n333_), .A4(new_n720_), .ZN(new_n751_));
  INV_X1    g550(.A(G50gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n725_), .B2(new_n431_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1331gat));
  NAND4_X1  g553(.A1(new_n635_), .A2(new_n680_), .A3(new_n681_), .A4(new_n444_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n442_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n669_), .A2(new_n505_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n678_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n679_), .A2(G57gat), .ZN(new_n759_));
  OAI22_X1  g558(.A1(new_n756_), .A2(G57gat), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT112), .ZN(G1332gat));
  OAI21_X1  g560(.A(G64gat), .B1(new_n758_), .B2(new_n732_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT48), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n732_), .A2(G64gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n755_), .B2(new_n764_), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n758_), .B2(new_n698_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT49), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n698_), .A2(G71gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n755_), .B2(new_n768_), .ZN(G1334gat));
  OAI21_X1  g568(.A(G78gat), .B1(new_n758_), .B2(new_n431_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT50), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n431_), .A2(G78gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n755_), .B2(new_n772_), .ZN(G1335gat));
  NOR3_X1   g572(.A1(new_n669_), .A2(new_n505_), .A3(new_n723_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n679_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n714_), .A2(new_n715_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n680_), .A2(new_n681_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(new_n677_), .A3(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n442_), .A2(new_n394_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1336gat));
  AOI21_X1  g579(.A(G92gat), .B1(new_n774_), .B2(new_n739_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n732_), .A2(new_n507_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n778_), .B2(new_n782_), .ZN(G1337gat));
  NAND3_X1  g582(.A1(new_n774_), .A2(new_n529_), .A3(new_n433_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n777_), .A2(new_n677_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n268_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n786_), .A2(KEYINPUT113), .A3(G99gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n786_), .B2(G99gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n774_), .A2(new_n524_), .A3(new_n333_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n785_), .B(new_n333_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G106gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n637_), .A2(new_n638_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n580_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n652_), .A2(new_n640_), .B1(new_n799_), .B2(new_n641_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n645_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n647_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n803_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n800_), .B(KEYINPUT55), .C1(new_n801_), .C2(new_n647_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n646_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n645_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n643_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n805_), .A2(new_n806_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n657_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT114), .B1(new_n650_), .B2(KEYINPUT55), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n807_), .A4(new_n810_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n658_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n813_), .A2(new_n661_), .A3(new_n505_), .A4(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n495_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n448_), .B1(new_n490_), .B2(new_n477_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n494_), .B1(new_n492_), .B2(new_n486_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n663_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n610_), .B1(new_n821_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT57), .B(new_n610_), .C1(new_n821_), .C2(new_n827_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n813_), .A2(new_n661_), .A3(new_n818_), .A4(new_n825_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT116), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT58), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(KEYINPUT116), .A3(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n834_), .A2(new_n611_), .A3(new_n613_), .A4(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n830_), .A2(new_n831_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n634_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n838_), .B2(new_n634_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n505_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n614_), .A2(new_n677_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n840_), .A2(new_n841_), .A3(new_n845_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n739_), .A2(new_n442_), .A3(new_n434_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT117), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT119), .B1(new_n846_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n838_), .A2(new_n634_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT118), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n843_), .B(KEYINPUT54), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n838_), .A2(new_n839_), .A3(new_n634_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  INV_X1    g656(.A(new_n850_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(new_n852_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n848_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT59), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n681_), .A2(new_n209_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n851_), .A2(new_n859_), .A3(new_n862_), .A4(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n209_), .B1(new_n861_), .B2(new_n681_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1340gat));
  INV_X1    g665(.A(new_n669_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n851_), .A2(new_n867_), .A3(new_n859_), .A4(new_n862_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G120gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n207_), .A2(KEYINPUT60), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n207_), .B1(new_n668_), .B2(KEYINPUT60), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n872_), .B2(new_n871_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n861_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n869_), .A2(new_n875_), .ZN(G1341gat));
  NOR2_X1   g675(.A1(new_n634_), .A2(new_n202_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n851_), .A2(new_n859_), .A3(new_n862_), .A4(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n202_), .B1(new_n861_), .B2(new_n634_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1342gat));
  NOR2_X1   g679(.A1(new_n614_), .A2(new_n203_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n851_), .A2(new_n859_), .A3(new_n862_), .A4(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n203_), .B1(new_n861_), .B2(new_n610_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1343gat));
  INV_X1    g683(.A(new_n430_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n860_), .A2(new_n885_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n886_), .A2(new_n442_), .A3(new_n731_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n505_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n867_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT121), .B(G148gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1345gat));
  NAND2_X1  g691(.A1(new_n887_), .A2(new_n677_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n887_), .B2(new_n722_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n614_), .A2(new_n305_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n887_), .B2(new_n897_), .ZN(G1347gat));
  XOR2_X1   g697(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n732_), .A2(new_n679_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(new_n698_), .A3(new_n333_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n856_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n681_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n900_), .B1(new_n905_), .B2(new_n236_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n246_), .ZN(new_n907_));
  OAI211_X1 g706(.A(G169gat), .B(new_n899_), .C1(new_n904_), .C2(new_n681_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1348gat));
  INV_X1    g708(.A(new_n904_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G176gat), .B1(new_n910_), .B2(new_n680_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n860_), .A2(new_n903_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n669_), .A2(new_n237_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n912_), .A2(KEYINPUT123), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT123), .B1(new_n912_), .B2(new_n913_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n911_), .A2(new_n914_), .A3(new_n915_), .ZN(G1349gat));
  AOI21_X1  g715(.A(G183gat), .B1(new_n912_), .B2(new_n677_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n634_), .A2(new_n230_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n910_), .B2(new_n918_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n904_), .B2(new_n614_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n722_), .A2(new_n231_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n904_), .B2(new_n921_), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n886_), .A2(new_n902_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n505_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g724(.A(new_n669_), .B1(KEYINPUT124), .B2(G204gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT125), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n927_), .B(new_n930_), .ZN(G1353gat));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n932_));
  INV_X1    g731(.A(G211gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n677_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT126), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n923_), .A2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n933_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1354gat));
  AND2_X1   g737(.A1(new_n615_), .A2(G218gat), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n860_), .A2(new_n885_), .A3(new_n901_), .A4(new_n939_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n886_), .A2(new_n610_), .A3(new_n902_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(G218gat), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT127), .B(new_n940_), .C1(new_n941_), .C2(G218gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1355gat));
endmodule


