//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NOR3_X1   g001(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT2), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n215_));
  OR3_X1    g014(.A1(new_n212_), .A2(new_n215_), .A3(KEYINPUT1), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n211_), .A4(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n206_), .A2(new_n208_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G127gat), .B(G134gat), .Z(new_n223_));
  XOR2_X1   g022(.A(G113gat), .B(G120gat), .Z(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT4), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n210_), .A2(new_n213_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n225_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(KEYINPUT4), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G1gat), .B(G29gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G85gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT0), .B(G57gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n226_), .A2(new_n230_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n233_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n235_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT91), .ZN(new_n243_));
  INV_X1    g042(.A(new_n239_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n233_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n241_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT19), .ZN(new_n250_));
  INV_X1    g049(.A(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n251_), .B2(G204gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n252_), .A2(new_n253_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT21), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G211gat), .B(G218gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n252_), .A2(KEYINPUT84), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(KEYINPUT84), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n259_), .B(new_n260_), .C1(new_n251_), .C2(G204gat), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n257_), .B(new_n258_), .C1(KEYINPUT21), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n262_), .A2(KEYINPUT86), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT86), .B1(new_n262_), .B2(new_n265_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G183gat), .ZN(new_n270_));
  INV_X1    g069(.A(G190gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT23), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT77), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT23), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT87), .Z(new_n281_));
  INV_X1    g080(.A(G176gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT24), .A3(new_n280_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(KEYINPUT24), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n275_), .A2(new_n272_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n279_), .A2(new_n284_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n267_), .A2(new_n269_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n262_), .A2(new_n265_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n276_), .A2(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n278_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G169gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT20), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n250_), .B1(new_n294_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n295_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(new_n293_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT20), .B1(new_n295_), .B2(new_n301_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n250_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT18), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT32), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n235_), .A2(KEYINPUT91), .A3(new_n239_), .A4(new_n241_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n250_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n305_), .A2(new_n293_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n250_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(KEYINPUT20), .A3(new_n320_), .A4(new_n302_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n314_), .A3(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n248_), .A2(new_n316_), .A3(new_n317_), .A4(new_n322_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT33), .B(new_n244_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT88), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT90), .B1(new_n232_), .B2(new_n234_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n239_), .B1(new_n240_), .B2(new_n233_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n328_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n227_), .A2(new_n331_), .A3(new_n233_), .A4(new_n231_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n326_), .A2(new_n329_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n318_), .A2(new_n313_), .A3(new_n321_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n313_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n247_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n323_), .B1(new_n325_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G233gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT82), .A2(G228gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(KEYINPUT82), .A2(G228gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n295_), .B(new_n346_), .C1(new_n347_), .C2(new_n228_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(KEYINPUT85), .A3(new_n295_), .A4(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n345_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G78gat), .B(G106gat), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n353_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n222_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G22gat), .B(G50gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n366_));
  OAI22_X1  g165(.A1(new_n358_), .A2(new_n359_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n353_), .A2(new_n355_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n356_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n365_), .A2(new_n366_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n353_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n340_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n367_), .A2(new_n372_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n248_), .A2(new_n317_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT27), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT92), .B(new_n379_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n313_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n309_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n334_), .A2(new_n379_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n382_), .A2(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n374_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G227gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(G15gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n394_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n296_), .A2(new_n399_), .A3(new_n300_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n301_), .A2(KEYINPUT30), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(KEYINPUT79), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT31), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n395_), .A2(new_n397_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT78), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(new_n400_), .A3(new_n401_), .A4(new_n398_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n404_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n229_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n403_), .A2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT31), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n225_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n382_), .A2(new_n383_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n385_), .A2(new_n386_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n373_), .A3(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n410_), .A2(new_n414_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n376_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT93), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n376_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n422_), .A2(new_n415_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n387_), .A4(new_n373_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n389_), .A2(new_n415_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT71), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT9), .ZN(new_n428_));
  INV_X1    g227(.A(G85gat), .ZN(new_n429_));
  INV_X1    g228(.A(G92gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G85gat), .A2(G92gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n428_), .B(new_n431_), .C1(new_n433_), .C2(KEYINPUT66), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n435_), .A2(KEYINPUT6), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(KEYINPUT6), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT10), .B(G99gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT65), .B(G106gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n431_), .A2(new_n442_), .A3(KEYINPUT9), .A4(new_n432_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n434_), .A2(new_n438_), .A3(new_n441_), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n445_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT7), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .A4(KEYINPUT67), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n446_), .B(new_n450_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT8), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n433_), .A2(KEYINPUT68), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n444_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G36gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G29gat), .ZN(new_n458_));
  INV_X1    g257(.A(G29gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G36gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G50gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G43gat), .ZN(new_n463_));
  INV_X1    g262(.A(G43gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G50gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n458_), .A2(new_n460_), .A3(new_n463_), .A4(new_n465_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT15), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n468_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n456_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n444_), .B(new_n470_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G232gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT34), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n477_), .A2(KEYINPUT35), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT69), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(KEYINPUT69), .A3(new_n478_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n477_), .A2(KEYINPUT35), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n474_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT70), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n473_), .A2(KEYINPUT70), .A3(new_n474_), .A4(new_n484_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n481_), .A2(new_n482_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G190gat), .B(G218gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G134gat), .B(G162gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT36), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n427_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n482_), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT69), .B1(new_n475_), .B2(new_n478_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n487_), .A2(new_n488_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT71), .B(new_n493_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n492_), .A2(KEYINPUT36), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n495_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n503_), .A2(KEYINPUT94), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(KEYINPUT94), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n426_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n511_));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n511_), .A2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n456_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n515_), .B(new_n444_), .C1(new_n455_), .C2(new_n454_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT12), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n456_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G230gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT64), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G120gat), .B(G148gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT5), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G176gat), .B(G204gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n517_), .A2(new_n518_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n525_), .B(new_n529_), .C1(new_n524_), .C2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n529_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n524_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n524_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT13), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G1gat), .A2(G8gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT14), .ZN(new_n541_));
  NOR2_X1   g340(.A1(G15gat), .A2(G22gat), .ZN(new_n542_));
  AND2_X1   g341(.A1(G15gat), .A2(G22gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G8gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n202_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n540_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n549_), .A2(new_n540_), .A3(new_n546_), .A4(new_n541_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n515_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555_));
  XOR2_X1   g354(.A(G127gat), .B(G155gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  OR3_X1    g358(.A1(new_n554_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(KEYINPUT17), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n544_), .A2(new_n547_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n549_), .A2(new_n541_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n468_), .B(new_n467_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n468_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n458_), .A2(new_n460_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n548_), .B(new_n550_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT74), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(new_n575_), .A3(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n472_), .A2(new_n469_), .A3(new_n551_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G169gat), .B(G197gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n575_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n586_));
  AOI211_X1 g385(.A(KEYINPUT74), .B(new_n571_), .C1(new_n566_), .C2(new_n569_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n579_), .B(new_n583_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n585_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n577_), .A2(KEYINPUT75), .A3(new_n579_), .A4(new_n583_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n588_), .A2(new_n589_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(KEYINPUT76), .A3(new_n585_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n539_), .A2(new_n563_), .A3(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n508_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n202_), .B1(new_n602_), .B2(new_n422_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT95), .Z(new_n604_));
  OAI21_X1  g403(.A(new_n502_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT37), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT72), .B(KEYINPUT37), .Z(new_n607_));
  NAND4_X1  g406(.A1(new_n495_), .A2(new_n500_), .A3(new_n502_), .A4(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n563_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n538_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT73), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n613_), .A2(new_n426_), .A3(new_n600_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n202_), .A3(new_n422_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n604_), .A2(new_n616_), .ZN(G1324gat));
  NAND2_X1  g416(.A1(new_n416_), .A2(new_n417_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n545_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n508_), .A2(new_n620_), .A3(new_n618_), .A4(new_n601_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(G8gat), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n508_), .A2(new_n618_), .A3(new_n601_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT96), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n622_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n623_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n619_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1325gat));
  AOI21_X1  g429(.A(new_n391_), .B1(new_n602_), .B2(new_n419_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n614_), .A2(new_n391_), .A3(new_n419_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n602_), .B2(new_n375_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT42), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n614_), .A2(new_n635_), .A3(new_n375_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1327gat));
  NOR2_X1   g438(.A1(new_n426_), .A2(new_n600_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n563_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n539_), .A2(new_n503_), .A3(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n459_), .A3(new_n422_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n538_), .A2(new_n563_), .A3(new_n599_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT97), .Z(new_n646_));
  OR2_X1    g445(.A1(new_n609_), .A2(KEYINPUT98), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT43), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n426_), .B2(new_n609_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n421_), .A2(new_n425_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n419_), .B1(new_n374_), .B2(new_n388_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n610_), .B(new_n648_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n646_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT44), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n653_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n646_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n654_), .A2(KEYINPUT99), .A3(KEYINPUT44), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n422_), .B(new_n655_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n663_), .A2(KEYINPUT100), .A3(G29gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT100), .B1(new_n663_), .B2(G29gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n644_), .B1(new_n664_), .B2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(KEYINPUT102), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n618_), .B(new_n655_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n667_), .A2(KEYINPUT102), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n387_), .A2(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n643_), .B2(new_n674_), .ZN(new_n675_));
  AND4_X1   g474(.A1(new_n640_), .A2(new_n642_), .A3(new_n673_), .A4(new_n674_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n669_), .B1(new_n671_), .B2(new_n678_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n668_), .B(new_n677_), .C1(new_n670_), .C2(G36gat), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  AOI21_X1  g480(.A(G43gat), .B1(new_n643_), .B2(new_n419_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n659_), .A2(new_n656_), .A3(new_n660_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT99), .B1(new_n654_), .B2(KEYINPUT44), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n683_), .A2(new_n684_), .B1(KEYINPUT44), .B2(new_n654_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n415_), .A2(new_n464_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT103), .B(KEYINPUT47), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1330gat));
  AOI21_X1  g488(.A(G50gat), .B1(new_n643_), .B2(new_n375_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n373_), .A2(new_n462_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n685_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n426_), .A2(new_n599_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(new_n539_), .A3(new_n611_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n422_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT104), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n599_), .A2(new_n563_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n508_), .A2(new_n539_), .A3(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT105), .B(G57gat), .Z(new_n699_));
  NOR2_X1   g498(.A1(new_n376_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n698_), .B2(new_n700_), .ZN(G1332gat));
  INV_X1    g500(.A(G64gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n698_), .B2(new_n618_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT48), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n694_), .A2(new_n702_), .A3(new_n618_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1333gat));
  INV_X1    g505(.A(G71gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n698_), .B2(new_n419_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n694_), .A2(new_n707_), .A3(new_n419_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1334gat));
  INV_X1    g511(.A(G78gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n698_), .B2(new_n375_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT50), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n694_), .A2(new_n713_), .A3(new_n375_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1335gat));
  AND3_X1   g516(.A1(new_n495_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n693_), .A2(new_n718_), .A3(new_n563_), .A4(new_n539_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT107), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n422_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n538_), .A2(new_n641_), .A3(new_n599_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n657_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(KEYINPUT108), .ZN(new_n724_));
  INV_X1    g523(.A(new_n722_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n724_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n376_), .A2(new_n429_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n721_), .B1(new_n729_), .B2(new_n730_), .ZN(G1336gat));
  NAND3_X1  g530(.A1(new_n720_), .A2(new_n430_), .A3(new_n618_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n724_), .A2(new_n387_), .A3(new_n728_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n430_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT109), .ZN(G1337gat));
  NAND3_X1  g534(.A1(new_n720_), .A2(new_n439_), .A3(new_n419_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G99gat), .B1(new_n723_), .B2(new_n415_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n720_), .A2(new_n440_), .A3(new_n375_), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT52), .B(new_n449_), .C1(new_n726_), .C2(new_n375_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n726_), .A2(new_n375_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G106gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n533_), .A2(KEYINPUT111), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(new_n751_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n525_), .B2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n522_), .A2(KEYINPUT55), .A3(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n532_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n750_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n522_), .A2(KEYINPUT55), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n761_), .B1(new_n534_), .B2(new_n755_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n529_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n762_), .A2(new_n748_), .A3(new_n763_), .A4(new_n749_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n599_), .A2(new_n531_), .A3(new_n760_), .A4(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n578_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n583_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n595_), .A2(new_n596_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n537_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n718_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n747_), .B(KEYINPUT57), .C1(new_n770_), .C2(KEYINPUT113), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n762_), .B(new_n763_), .C1(KEYINPUT114), .C2(KEYINPUT56), .ZN(new_n772_));
  NOR2_X1   g571(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n531_), .A2(new_n768_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n777_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n610_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n597_), .A2(KEYINPUT76), .A3(new_n585_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT76), .B1(new_n597_), .B2(new_n585_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n531_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n760_), .A2(new_n764_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n769_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n503_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT115), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n788_), .B2(KEYINPUT115), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n771_), .B(new_n782_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n563_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n697_), .A2(KEYINPUT110), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n697_), .A2(KEYINPUT110), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n795_), .A2(new_n538_), .A3(new_n609_), .A4(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT54), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n794_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n418_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n415_), .A2(new_n376_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n803_));
  INV_X1    g602(.A(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n793_), .A2(new_n806_), .A3(new_n563_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NOR4_X1   g607(.A1(new_n418_), .A2(KEYINPUT59), .A3(new_n376_), .A4(new_n415_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n803_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT117), .B(G113gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n599_), .A2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT118), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n802_), .A2(new_n600_), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n811_), .A2(new_n814_), .B1(G113gat), .B2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT119), .ZN(G1340gat));
  OAI21_X1  g616(.A(G120gat), .B1(new_n811_), .B2(new_n538_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n802_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n820_));
  AOI21_X1  g619(.A(G120gat), .B1(new_n539_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n820_), .B2(G120gat), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n819_), .B(new_n822_), .C1(new_n821_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n818_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT121), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n818_), .A2(new_n828_), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1341gat));
  OAI21_X1  g629(.A(G127gat), .B1(new_n811_), .B2(new_n563_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n563_), .A2(G127gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n802_), .B2(new_n832_), .ZN(G1342gat));
  OAI21_X1  g632(.A(G134gat), .B1(new_n811_), .B2(new_n609_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n802_), .A2(G134gat), .A3(new_n506_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(KEYINPUT122), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1343gat));
  NOR4_X1   g639(.A1(new_n618_), .A2(new_n373_), .A3(new_n419_), .A4(new_n376_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n799_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n599_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n539_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g646(.A1(new_n842_), .A2(new_n563_), .ZN(new_n848_));
  XOR2_X1   g647(.A(KEYINPUT61), .B(G155gat), .Z(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  OAI21_X1  g649(.A(G162gat), .B1(new_n842_), .B2(new_n609_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n506_), .A2(G162gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n842_), .B2(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n420_), .A2(new_n387_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n373_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n808_), .B2(new_n856_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n793_), .A2(new_n806_), .A3(new_n563_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n806_), .B1(new_n793_), .B2(new_n563_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n798_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n856_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT124), .A3(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n857_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n283_), .A3(new_n599_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n855_), .A2(new_n599_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT123), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n373_), .ZN(new_n867_));
  OAI21_X1  g666(.A(G169gat), .B1(new_n808_), .B2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT62), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n869_), .ZN(G1348gat));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  INV_X1    g670(.A(new_n799_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n375_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n799_), .A2(KEYINPUT125), .A3(new_n373_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n855_), .A3(new_n874_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n875_), .A2(new_n282_), .A3(new_n538_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n863_), .A2(new_n539_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n282_), .ZN(G1349gat));
  OR2_X1    g677(.A1(new_n875_), .A2(new_n563_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n563_), .A2(new_n285_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n879_), .A2(new_n270_), .B1(new_n863_), .B2(new_n880_), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n857_), .A2(new_n610_), .A3(new_n862_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G190gat), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n857_), .A2(new_n507_), .A3(new_n286_), .A4(new_n862_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT126), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(new_n887_), .A3(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1351gat));
  NAND3_X1  g688(.A1(new_n378_), .A2(new_n618_), .A3(new_n415_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n872_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n600_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n251_), .A2(KEYINPUT127), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n251_), .A2(KEYINPUT127), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n893_), .B2(new_n895_), .ZN(G1352gat));
  NAND2_X1  g696(.A1(new_n891_), .A2(new_n539_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g698(.A1(new_n891_), .A2(new_n641_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  OR3_X1    g703(.A1(new_n892_), .A2(G218gat), .A3(new_n506_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G218gat), .B1(new_n892_), .B2(new_n609_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1355gat));
endmodule


