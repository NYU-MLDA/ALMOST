//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(G134gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT78), .B(G127gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n207_), .A3(new_n205_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT79), .Z(new_n212_));
  INV_X1    g011(.A(KEYINPUT31), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT23), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT22), .B(G169gat), .Z(new_n219_));
  OAI211_X1 g018(.A(new_n217_), .B(new_n218_), .C1(G176gat), .C2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(KEYINPUT26), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n223_), .B(new_n224_), .C1(new_n225_), .C2(new_n221_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n227_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n226_), .A2(new_n216_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n220_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G43gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT30), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n233_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G15gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  AND3_X1   g042(.A1(new_n235_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n214_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT81), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n239_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n243_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n212_), .B(KEYINPUT31), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n235_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT80), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT3), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT2), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n263_), .A2(new_n266_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n260_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n257_), .A2(KEYINPUT1), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT82), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT82), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n257_), .A2(new_n274_), .A3(KEYINPUT1), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n275_), .A3(new_n256_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n257_), .A2(KEYINPUT1), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n264_), .B(new_n262_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(G197gat), .B(G204gat), .Z(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G106gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G228gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(G78gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G106gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n280_), .A2(new_n291_), .A3(new_n285_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n287_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n287_), .B2(new_n292_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT84), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n287_), .A2(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n290_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n287_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G22gat), .B(G50gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n302_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n302_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n305_), .A3(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n295_), .A2(new_n301_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n311_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n314_), .A2(new_n299_), .A3(new_n300_), .A4(new_n298_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n255_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT27), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n283_), .B(new_n284_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n220_), .A3(new_n232_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n225_), .A2(new_n224_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n216_), .A2(KEYINPUT85), .A3(new_n229_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT85), .B1(new_n216_), .B2(new_n229_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n231_), .B(new_n321_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n220_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n285_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n325_), .B2(new_n285_), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT20), .B(new_n320_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT89), .ZN(new_n334_));
  XOR2_X1   g133(.A(G64gat), .B(G92gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n319_), .A2(new_n324_), .A3(new_n220_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n331_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n285_), .A2(new_n233_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT20), .A4(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n332_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n339_), .B1(new_n332_), .B2(new_n345_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n318_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT99), .ZN(new_n349_));
  INV_X1    g148(.A(new_n331_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT20), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n325_), .A2(new_n285_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT86), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n325_), .A2(new_n326_), .A3(new_n285_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n355_), .B2(new_n320_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n345_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n338_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n332_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT99), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n318_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n349_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT98), .B1(new_n329_), .B2(new_n331_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT98), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n355_), .A2(new_n365_), .A3(new_n350_), .A4(new_n320_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n367_));
  AND3_X1   g166(.A1(new_n344_), .A2(new_n340_), .A3(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n364_), .B(new_n366_), .C1(new_n350_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n338_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(KEYINPUT27), .A3(new_n359_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n363_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT93), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n375_));
  NAND3_X1  g174(.A1(new_n211_), .A2(new_n279_), .A3(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n271_), .A2(new_n278_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n210_), .A4(new_n209_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT92), .B1(new_n211_), .B2(new_n279_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n211_), .A2(new_n279_), .A3(KEYINPUT91), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT91), .B1(new_n211_), .B2(new_n279_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n379_), .B(new_n380_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n374_), .B(new_n376_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n383_), .A2(new_n374_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n385_), .A2(new_n386_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n317_), .A2(new_n372_), .A3(new_n396_), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n393_), .A2(new_n313_), .A3(new_n395_), .A4(new_n315_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n361_), .B1(new_n360_), .B2(new_n318_), .ZN(new_n399_));
  AOI211_X1 g198(.A(KEYINPUT99), .B(KEYINPUT27), .C1(new_n358_), .C2(new_n359_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n398_), .B(new_n371_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT100), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n339_), .A2(KEYINPUT32), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n332_), .A2(new_n404_), .A3(new_n345_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n332_), .A2(new_n404_), .A3(KEYINPUT96), .A4(new_n345_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n404_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n369_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n396_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n395_), .A2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n381_), .A2(new_n382_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n374_), .A3(new_n380_), .A4(new_n379_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n376_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n392_), .B(new_n416_), .C1(new_n417_), .C2(new_n374_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n395_), .A2(new_n413_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT90), .B1(new_n346_), .B2(new_n347_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n358_), .A2(new_n422_), .A3(new_n359_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n412_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n316_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n363_), .A2(KEYINPUT100), .A3(new_n398_), .A4(new_n371_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n403_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n255_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n397_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT70), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G232gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT34), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT66), .B(KEYINPUT35), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT69), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT7), .ZN(new_n437_));
  INV_X1    g236(.A(G99gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n291_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n438_), .A2(KEYINPUT10), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n438_), .A2(KEYINPUT10), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n291_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n442_), .A2(new_n443_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(KEYINPUT9), .A3(new_n447_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n447_), .A2(KEYINPUT9), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .A4(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n445_), .A2(KEYINPUT8), .A3(new_n448_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n238_), .A2(G50gat), .ZN(new_n461_));
  INV_X1    g260(.A(G50gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(G43gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G29gat), .A2(G36gat), .ZN(new_n464_));
  AND2_X1   g263(.A1(G29gat), .A2(G36gat), .ZN(new_n465_));
  OAI22_X1  g264(.A1(new_n461_), .A2(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n462_), .A2(G43gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n238_), .A2(G50gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G29gat), .A2(G36gat), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n471_), .A3(KEYINPUT15), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n436_), .B1(new_n460_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n472_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n451_), .A2(new_n479_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n433_), .A2(new_n434_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n435_), .A2(KEYINPUT69), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n431_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n480_), .A2(new_n481_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n485_), .A2(new_n477_), .A3(KEYINPUT70), .A4(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n460_), .A2(new_n476_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT67), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n460_), .A2(new_n489_), .A3(new_n476_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n484_), .A2(new_n486_), .B1(new_n491_), .B2(new_n435_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G190gat), .B(G218gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G134gat), .B(G162gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(KEYINPUT36), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n497_), .A2(KEYINPUT36), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n492_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n492_), .B2(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n430_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(KEYINPUT71), .A2(G22gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G15gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(KEYINPUT71), .A2(G22gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(KEYINPUT71), .A2(G22gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(G15gat), .B1(new_n510_), .B2(new_n505_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(G1gat), .B2(G8gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G8gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n517_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n519_), .A3(new_n515_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(G231gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(G57gat), .A2(G64gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G57gat), .A2(G64gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT11), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G71gat), .B(G78gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT11), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n530_), .A3(new_n525_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n528_), .A3(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n523_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n523_), .A2(new_n534_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT73), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT16), .B(G183gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT17), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(KEYINPUT17), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n538_), .A2(new_n541_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n546_), .B(KEYINPUT72), .Z(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT65), .ZN(new_n552_));
  XOR2_X1   g351(.A(G176gat), .B(G204gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT64), .B(KEYINPUT5), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n532_), .A2(new_n533_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n460_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n534_), .A2(new_n451_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(KEYINPUT12), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n460_), .A2(new_n562_), .A3(new_n558_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n565_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n557_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n565_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n557_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n571_), .A2(new_n567_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n552_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n568_), .A3(new_n557_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n572_), .B1(new_n571_), .B2(new_n567_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(KEYINPUT65), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n519_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n514_), .B(new_n517_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n466_), .A2(new_n471_), .A3(KEYINPUT15), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT15), .B1(new_n466_), .B2(new_n471_), .ZN(new_n584_));
  OAI22_X1  g383(.A1(new_n581_), .A2(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT75), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n476_), .B(new_n587_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n518_), .A2(new_n520_), .A3(new_n479_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT76), .Z(new_n591_));
  NAND4_X1  g390(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .A4(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n479_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n581_), .A2(new_n582_), .A3(new_n472_), .ZN(new_n594_));
  OAI211_X1 g393(.A(G229gat), .B(G233gat), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n592_), .A2(new_n595_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n580_), .A2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n504_), .A2(new_n551_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n202_), .B1(new_n606_), .B2(new_n396_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT102), .Z(new_n608_));
  NAND2_X1  g407(.A1(new_n503_), .A2(KEYINPUT37), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n498_), .B(new_n610_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n609_), .A2(new_n551_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT74), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n430_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(new_n605_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n396_), .B(KEYINPUT101), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n202_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(G8gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(new_n620_), .A3(new_n372_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n606_), .A2(new_n372_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(G8gat), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n621_), .B(KEYINPUT40), .C1(new_n624_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  AOI21_X1  g429(.A(new_n507_), .B1(new_n606_), .B2(new_n255_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n615_), .A2(new_n507_), .A3(new_n255_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n316_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n615_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n606_), .B2(new_n636_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(G1327gat));
  INV_X1    g441(.A(new_n503_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n551_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n605_), .A2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n430_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n396_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n645_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n428_), .A2(new_n429_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n397_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n609_), .A2(new_n611_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n430_), .A2(KEYINPUT43), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n648_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT44), .B(new_n648_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n616_), .A2(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n647_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  XNOR2_X1  g462(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(new_n372_), .A3(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G36gat), .ZN(new_n666_));
  INV_X1    g465(.A(G36gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n646_), .A2(new_n667_), .A3(new_n372_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT45), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n646_), .A2(KEYINPUT45), .A3(new_n667_), .A4(new_n372_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n664_), .B1(new_n666_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n664_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n672_), .B(new_n675_), .C1(new_n665_), .C2(G36gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1329gat));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n659_), .A2(new_n255_), .A3(new_n660_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G43gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n646_), .A2(new_n238_), .A3(new_n255_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n681_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT47), .B(new_n683_), .C1(new_n679_), .C2(G43gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1330gat));
  NAND3_X1  g484(.A1(new_n659_), .A2(new_n636_), .A3(new_n660_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT106), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n659_), .A2(new_n688_), .A3(new_n636_), .A4(new_n660_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(G50gat), .A3(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n646_), .A2(new_n462_), .A3(new_n636_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1331gat));
  XNOR2_X1  g491(.A(new_n578_), .B(KEYINPUT13), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n603_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n614_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G57gat), .B1(new_n695_), .B2(new_n616_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n504_), .A2(new_n551_), .A3(new_n694_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n396_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT107), .B(G57gat), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(G1332gat));
  INV_X1    g500(.A(G64gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n695_), .A2(new_n702_), .A3(new_n372_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n372_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G64gat), .B1(new_n697_), .B2(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT108), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(KEYINPUT108), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n703_), .B1(new_n709_), .B2(new_n710_), .ZN(G1333gat));
  INV_X1    g510(.A(G71gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n695_), .A2(new_n712_), .A3(new_n255_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n697_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n714_), .B2(new_n255_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n716_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n697_), .B2(new_n316_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n695_), .A2(new_n289_), .A3(new_n636_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n694_), .A2(new_n644_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n430_), .A2(new_n643_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n616_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n654_), .A2(new_n656_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n724_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n396_), .A2(G85gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n725_), .B2(new_n372_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT110), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n372_), .A2(G92gat), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT111), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n728_), .B2(new_n734_), .ZN(G1337gat));
  OAI211_X1 g534(.A(new_n725_), .B(new_n255_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n727_), .A2(new_n429_), .A3(new_n724_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n438_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n725_), .A2(new_n291_), .A3(new_n636_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n724_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n636_), .B(new_n741_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(G106gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G106gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n740_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n740_), .B(new_n747_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1339gat));
  INV_X1    g550(.A(new_n591_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .A4(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n591_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n599_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT115), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n753_), .A2(new_n754_), .A3(new_n757_), .A4(new_n599_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n602_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n575_), .A2(KEYINPUT65), .A3(new_n576_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT65), .B1(new_n575_), .B2(new_n576_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n578_), .A2(KEYINPUT116), .A3(new_n760_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n564_), .A2(KEYINPUT55), .A3(new_n565_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n561_), .A2(new_n570_), .A3(new_n563_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n770_));
  NOR2_X1   g569(.A1(new_n571_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT56), .B(new_n572_), .C1(new_n769_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n767_), .B(new_n768_), .C1(new_n571_), .C2(new_n770_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n572_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n603_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n572_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(KEYINPUT114), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n575_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n765_), .B(new_n766_), .C1(new_n777_), .C2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(KEYINPUT57), .A3(new_n643_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT118), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n643_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n778_), .A2(new_n779_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(KEYINPUT117), .A3(new_n772_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n775_), .A2(new_n790_), .A3(KEYINPUT56), .A4(new_n572_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(new_n575_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n792_), .A3(new_n760_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n789_), .A2(new_n792_), .A3(KEYINPUT58), .A4(new_n760_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n653_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n782_), .A2(new_n798_), .A3(KEYINPUT57), .A4(new_n643_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n784_), .A2(new_n787_), .A3(new_n797_), .A4(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n644_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n612_), .A2(new_n802_), .A3(new_n604_), .A4(new_n693_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n609_), .A2(new_n551_), .A3(new_n604_), .A4(new_n611_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT54), .B1(new_n804_), .B2(new_n580_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT119), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n809_), .B(new_n806_), .C1(new_n800_), .C2(new_n644_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n704_), .A2(new_n616_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n811_), .A2(new_n317_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n808_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT120), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT116), .B1(new_n578_), .B2(new_n760_), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n764_), .B(new_n759_), .C1(new_n574_), .C2(new_n577_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n788_), .A2(new_n773_), .A3(new_n772_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(new_n603_), .A3(new_n575_), .A4(new_n780_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n503_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n798_), .B1(new_n820_), .B2(KEYINPUT57), .ZN(new_n821_));
  INV_X1    g620(.A(new_n799_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n795_), .A2(new_n796_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n824_), .A2(new_n653_), .B1(new_n786_), .B2(new_n785_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n551_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n809_), .B1(new_n826_), .B2(new_n806_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n801_), .A2(KEYINPUT119), .A3(new_n807_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n811_), .A2(new_n317_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n827_), .A2(KEYINPUT120), .A3(new_n828_), .A4(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n603_), .B1(new_n814_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G113gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n826_), .A2(new_n806_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n812_), .A2(KEYINPUT121), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(KEYINPUT59), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n604_), .A2(new_n833_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n832_), .A2(new_n833_), .B1(new_n842_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(G120gat), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT60), .B1(new_n580_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n849_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n846_), .B(new_n848_), .C1(new_n850_), .C2(new_n830_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n842_), .B2(new_n580_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n813_), .A2(new_n836_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G120gat), .B1(new_n854_), .B2(new_n693_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n846_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n848_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n856_), .B(new_n857_), .C1(new_n814_), .C2(new_n831_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n855_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(new_n860_), .ZN(G1341gat));
  OAI21_X1  g660(.A(new_n551_), .B1(new_n814_), .B2(new_n831_), .ZN(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(KEYINPUT123), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n644_), .B1(new_n850_), .B2(new_n830_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(G127gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n644_), .A2(new_n863_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n864_), .A2(new_n867_), .B1(new_n842_), .B2(new_n868_), .ZN(G1342gat));
  OAI21_X1  g668(.A(new_n503_), .B1(new_n814_), .B2(new_n831_), .ZN(new_n870_));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n655_), .A2(new_n871_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n871_), .B1(new_n842_), .B2(new_n872_), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  INV_X1    g673(.A(new_n811_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n827_), .A2(new_n429_), .A3(new_n828_), .A4(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n876_), .B2(new_n316_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n808_), .A2(new_n810_), .A3(new_n255_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n878_), .A2(KEYINPUT124), .A3(new_n636_), .A4(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n603_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G141gat), .ZN(new_n882_));
  INV_X1    g681(.A(G141gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n883_), .A3(new_n603_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1344gat));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n580_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G148gat), .ZN(new_n887_));
  INV_X1    g686(.A(G148gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n880_), .A2(new_n888_), .A3(new_n580_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1345gat));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n880_), .B2(new_n551_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n891_), .ZN(new_n893_));
  AOI211_X1 g692(.A(new_n644_), .B(new_n893_), .C1(new_n877_), .C2(new_n879_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n880_), .B2(new_n503_), .ZN(new_n896_));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  AOI211_X1 g696(.A(new_n897_), .B(new_n655_), .C1(new_n877_), .C2(new_n879_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(G169gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n704_), .A2(new_n317_), .A3(new_n616_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n834_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n903_), .B2(new_n603_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n834_), .A2(new_n219_), .A3(new_n604_), .A4(new_n902_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT62), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(KEYINPUT62), .B2(new_n904_), .ZN(G1348gat));
  AOI21_X1  g706(.A(G176gat), .B1(new_n903_), .B2(new_n580_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n808_), .A2(new_n810_), .A3(new_n902_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n580_), .A2(G176gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1349gat));
  NOR4_X1   g710(.A1(new_n834_), .A2(new_n644_), .A3(new_n224_), .A4(new_n902_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n909_), .A2(new_n551_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(G183gat), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(KEYINPUT125), .B(new_n913_), .C1(new_n914_), .C2(G183gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1350gat));
  AOI21_X1  g718(.A(new_n222_), .B1(new_n903_), .B2(new_n653_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT126), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n903_), .A2(new_n225_), .A3(new_n503_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1351gat));
  NOR2_X1   g722(.A1(new_n808_), .A2(new_n810_), .ZN(new_n924_));
  AND4_X1   g723(.A1(new_n429_), .A2(new_n924_), .A3(new_n398_), .A4(new_n372_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n603_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n580_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n925_), .B2(new_n551_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n878_), .A2(new_n398_), .A3(new_n372_), .ZN(new_n932_));
  XOR2_X1   g731(.A(KEYINPUT63), .B(G211gat), .Z(new_n933_));
  NOR3_X1   g732(.A1(new_n932_), .A2(new_n644_), .A3(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT127), .B1(new_n931_), .B2(new_n934_), .ZN(new_n935_));
  OAI22_X1  g734(.A1(new_n932_), .A2(new_n644_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n925_), .A2(new_n551_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n936_), .B(new_n937_), .C1(new_n938_), .C2(new_n933_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n935_), .A2(new_n939_), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n925_), .B2(new_n503_), .ZN(new_n941_));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n932_), .A2(new_n942_), .A3(new_n655_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1355gat));
endmodule


