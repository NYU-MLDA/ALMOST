//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT73), .ZN(new_n203_));
  XOR2_X1   g002(.A(G127gat), .B(G155gat), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT17), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G1gat), .A2(G8gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT14), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G231gat), .A2(G233gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G57gat), .B(G64gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n219_));
  XOR2_X1   g018(.A(G71gat), .B(G78gat), .Z(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n220_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n218_), .A2(KEYINPUT11), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n217_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n207_), .A2(new_n208_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n209_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT75), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n209_), .A2(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT74), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT37), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G190gat), .B(G218gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G134gat), .B(G162gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT36), .Z(new_n236_));
  NAND2_X1  g035(.A1(G232gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT34), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT35), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT68), .Z(new_n240_));
  INV_X1    g039(.A(G85gat), .ZN(new_n241_));
  INV_X1    g040(.A(G92gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT6), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT6), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  INV_X1    g051(.A(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  OAI22_X1  g054(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n245_), .B1(new_n250_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT8), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT9), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n244_), .A2(new_n262_), .A3(new_n261_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n244_), .B2(new_n261_), .ZN(new_n264_));
  OAI221_X1 g063(.A(new_n243_), .B1(new_n261_), .B2(new_n244_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT10), .B(G99gat), .Z(new_n266_));
  AOI22_X1  g065(.A1(new_n266_), .A2(new_n254_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(KEYINPUT8), .B(new_n245_), .C1(new_n250_), .C2(new_n257_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G29gat), .B(G36gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G43gat), .B(G50gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OAI22_X1  g073(.A1(new_n270_), .A2(new_n274_), .B1(KEYINPUT35), .B2(new_n238_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(KEYINPUT67), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n273_), .B(KEYINPUT15), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n260_), .A2(new_n268_), .A3(new_n278_), .A4(new_n269_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n275_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n276_), .A2(KEYINPUT69), .A3(new_n277_), .A4(new_n279_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n240_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n240_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT70), .ZN(new_n286_));
  INV_X1    g085(.A(new_n275_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(KEYINPUT70), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n286_), .A2(new_n280_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n236_), .B1(new_n284_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n232_), .B1(new_n291_), .B2(KEYINPUT71), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n235_), .A2(KEYINPUT36), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n282_), .A2(new_n283_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n289_), .B(new_n293_), .C1(new_n294_), .C2(new_n240_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n295_), .B(new_n291_), .C1(KEYINPUT71), .C2(new_n232_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n231_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G230gat), .A2(G233gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n270_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n304_), .A2(new_n224_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n224_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n276_), .A2(new_n279_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT12), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n224_), .A2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n304_), .B2(new_n224_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n304_), .A2(new_n224_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n313_), .A2(new_n302_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT5), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G176gat), .B(G204gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n309_), .A2(new_n316_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT13), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(KEYINPUT13), .A3(new_n324_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n301_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT76), .ZN(new_n331_));
  XOR2_X1   g130(.A(G8gat), .B(G36gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT86), .ZN(new_n339_));
  INV_X1    g138(.A(G204gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(G197gat), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n340_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(G197gat), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(G197gat), .B2(G204gat), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n351_), .A2(KEYINPUT85), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT85), .B1(new_n351_), .B2(new_n353_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n338_), .B(new_n350_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n352_), .B(new_n338_), .C1(new_n344_), .C2(new_n348_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT22), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT22), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(G169gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n363_), .A3(KEYINPUT91), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT91), .B1(new_n361_), .B2(new_n363_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n365_), .A2(new_n366_), .A3(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT23), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G183gat), .ZN(new_n373_));
  INV_X1    g172(.A(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(KEYINPUT25), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G183gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n374_), .A2(KEYINPUT26), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT26), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G190gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT24), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n387_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT80), .B1(new_n369_), .B2(new_n371_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n368_), .B2(KEYINPUT23), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  OAI22_X1  g197(.A1(new_n367_), .A2(new_n380_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n337_), .B1(new_n359_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT94), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n338_), .ZN(new_n403_));
  AND2_X1   g202(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n406_), .A2(G197gat), .B1(new_n341_), .B2(new_n343_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n403_), .B1(new_n407_), .B2(new_n349_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n404_), .A2(new_n405_), .A3(G197gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT21), .B1(new_n342_), .B2(new_n340_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n351_), .A2(KEYINPUT85), .A3(new_n353_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n357_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n379_), .A2(KEYINPUT24), .A3(new_n389_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n387_), .A2(new_n372_), .A3(new_n393_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n375_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n418_));
  INV_X1    g217(.A(G176gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n361_), .A2(new_n363_), .A3(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n379_), .A2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n416_), .A2(new_n417_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT92), .B1(new_n415_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT92), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n416_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n418_), .A2(new_n421_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n359_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT94), .B(new_n337_), .C1(new_n359_), .C2(new_n399_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n402_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT19), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n431_), .A2(KEYINPUT95), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n359_), .B2(new_n399_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n433_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n415_), .A2(new_n422_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n431_), .A2(new_n433_), .B1(KEYINPUT95), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n336_), .B1(new_n434_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT96), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT96), .B(new_n336_), .C1(new_n434_), .C2(new_n440_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n433_), .A2(new_n435_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n359_), .B2(new_n399_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n429_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n366_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n419_), .A3(new_n364_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n380_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n398_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n394_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n450_), .A2(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT20), .B1(new_n454_), .B2(new_n415_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n359_), .A2(new_n427_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n433_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n448_), .A2(new_n335_), .A3(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(KEYINPUT27), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n443_), .A2(new_n444_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G155gat), .ZN(new_n461_));
  INV_X1    g260(.A(G162gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT1), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT82), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT82), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(G155gat), .B2(G162gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT1), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(G155gat), .A3(G162gat), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n463_), .A2(new_n464_), .A3(new_n466_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G141gat), .ZN(new_n470_));
  INV_X1    g269(.A(G148gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G141gat), .A2(G148gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT2), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT83), .B1(new_n472_), .B2(KEYINPUT3), .ZN(new_n481_));
  NOR3_X1   g280(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT83), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n480_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n464_), .B(new_n466_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n475_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G127gat), .B(G134gat), .Z(new_n488_));
  XOR2_X1   g287(.A(G113gat), .B(G120gat), .Z(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT4), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n481_), .A2(new_n484_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n480_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n486_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n475_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n488_), .B(new_n489_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n491_), .A3(KEYINPUT4), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G1gat), .B(G29gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G85gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT0), .B(G57gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n503_), .B1(new_n499_), .B2(new_n491_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n502_), .B1(new_n492_), .B2(new_n500_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n508_), .B1(new_n513_), .B2(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n422_), .B(KEYINPUT30), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G227gat), .A2(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(G15gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G71gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(new_n253_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n516_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n498_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n516_), .B(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n490_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT81), .B(G43gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT31), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n515_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n446_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n336_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT27), .B1(new_n536_), .B2(new_n458_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n497_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT28), .B1(new_n487_), .B2(KEYINPUT29), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G22gat), .B(G50gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n487_), .A2(KEYINPUT29), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n359_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G228gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n550_), .B(new_n552_), .C1(new_n553_), .C2(new_n415_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n359_), .B(new_n549_), .C1(KEYINPUT88), .C2(new_n551_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G78gat), .B(G106gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT90), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n548_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n415_), .B2(new_n553_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n356_), .A2(new_n358_), .B1(new_n487_), .B2(KEYINPUT29), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n555_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n556_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(KEYINPUT89), .B(new_n556_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n554_), .A2(KEYINPUT90), .A3(new_n555_), .A4(new_n557_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n560_), .A2(new_n567_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n558_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n548_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n460_), .A2(new_n533_), .A3(new_n538_), .A4(new_n573_), .ZN(new_n574_));
  AOI211_X1 g373(.A(new_n515_), .B(new_n537_), .C1(new_n570_), .C2(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n431_), .A2(new_n433_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n439_), .A2(KEYINPUT95), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n431_), .A2(KEYINPUT95), .A3(new_n433_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n576_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n448_), .A2(new_n457_), .A3(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n515_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n514_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT33), .B(new_n508_), .C1(new_n513_), .C2(new_n510_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n499_), .A2(new_n491_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n508_), .B1(new_n588_), .B2(new_n503_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n536_), .A3(new_n458_), .ZN(new_n591_));
  OAI22_X1  g390(.A1(new_n581_), .A2(new_n583_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n460_), .A2(new_n575_), .B1(new_n592_), .B2(new_n573_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n531_), .A2(new_n532_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n574_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n215_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n273_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n215_), .A2(new_n274_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n597_), .A2(KEYINPUT77), .A3(new_n598_), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n596_), .A2(KEYINPUT77), .A3(new_n273_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT78), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n277_), .A2(new_n215_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n601_), .A3(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G169gat), .B(G197gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  XOR2_X1   g409(.A(new_n607_), .B(new_n610_), .Z(new_n611_));
  AND2_X1   g410(.A1(new_n595_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n331_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT97), .ZN(new_n614_));
  INV_X1    g413(.A(new_n515_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(G1gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(KEYINPUT38), .A3(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n228_), .A2(new_n230_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n329_), .A2(new_n611_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT98), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n595_), .A2(new_n296_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n615_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT38), .B1(new_n614_), .B2(new_n616_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT99), .B(KEYINPUT38), .C1(new_n614_), .C2(new_n616_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n617_), .B(new_n623_), .C1(new_n626_), .C2(new_n627_), .ZN(G1324gat));
  NAND2_X1  g427(.A1(new_n460_), .A2(new_n538_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(G8gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n614_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n622_), .B2(new_n630_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n632_), .B(new_n637_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  NAND3_X1  g440(.A1(new_n620_), .A2(new_n594_), .A3(new_n621_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n642_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(new_n642_), .B2(G15gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n594_), .A2(new_n518_), .ZN(new_n645_));
  OAI22_X1  g444(.A1(new_n643_), .A2(new_n644_), .B1(new_n613_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT101), .ZN(G1326gat));
  OAI21_X1  g446(.A(G22gat), .B1(new_n622_), .B2(new_n573_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n573_), .A2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n613_), .B2(new_n650_), .ZN(G1327gat));
  INV_X1    g450(.A(new_n329_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n652_), .A2(new_n296_), .A3(new_n618_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n653_), .A2(new_n612_), .ZN(new_n654_));
  INV_X1    g453(.A(G29gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n515_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n595_), .A2(new_n658_), .A3(new_n300_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n460_), .A2(new_n575_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n592_), .A2(new_n573_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n594_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AND4_X1   g461(.A1(new_n460_), .A2(new_n533_), .A3(new_n538_), .A4(new_n573_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT102), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(new_n574_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n297_), .A2(KEYINPUT103), .A3(new_n298_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT103), .B1(new_n297_), .B2(new_n298_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(new_n666_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n659_), .B1(new_n671_), .B2(KEYINPUT43), .ZN(new_n672_));
  INV_X1    g471(.A(new_n611_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n652_), .A2(new_n673_), .A3(new_n618_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n657_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT104), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n657_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n669_), .B1(new_n595_), .B2(KEYINPUT102), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n658_), .B1(new_n680_), .B2(new_n666_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n674_), .C1(new_n681_), .C2(new_n659_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT105), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n671_), .A2(KEYINPUT43), .ZN(new_n684_));
  INV_X1    g483(.A(new_n659_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(KEYINPUT44), .A4(new_n674_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n677_), .A2(new_n679_), .B1(new_n683_), .B2(new_n688_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT106), .B(new_n655_), .C1(new_n689_), .C2(new_n515_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n677_), .A2(new_n679_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n683_), .A2(new_n688_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n515_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n691_), .B1(new_n694_), .B2(G29gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n656_), .B1(new_n690_), .B2(new_n695_), .ZN(G1328gat));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n689_), .B2(new_n629_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n654_), .A2(new_n698_), .A3(new_n629_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT45), .Z(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n692_), .A2(new_n629_), .A3(new_n693_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  INV_X1    g503(.A(new_n701_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(KEYINPUT46), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n706_), .ZN(G1329gat));
  NAND4_X1  g506(.A1(new_n692_), .A2(G43gat), .A3(new_n693_), .A4(new_n594_), .ZN(new_n708_));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n654_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n594_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  INV_X1    g516(.A(new_n573_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G50gat), .B1(new_n654_), .B2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(G50gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n689_), .B2(new_n720_), .ZN(G1331gat));
  AND2_X1   g520(.A1(new_n595_), .A2(new_n673_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n301_), .A3(new_n652_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT108), .ZN(new_n724_));
  INV_X1    g523(.A(G57gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(new_n515_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n329_), .A2(new_n231_), .A3(new_n611_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n621_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n615_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(new_n730_), .ZN(G1332gat));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n728_), .B2(new_n629_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT48), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n724_), .A2(new_n732_), .A3(new_n629_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n728_), .B2(new_n594_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT49), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n724_), .A2(new_n737_), .A3(new_n594_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n728_), .B2(new_n718_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT109), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT50), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(KEYINPUT50), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n724_), .A2(new_n742_), .A3(new_n718_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(G1335gat));
  OR2_X1    g547(.A1(new_n672_), .A2(KEYINPUT111), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n329_), .A2(new_n611_), .A3(new_n618_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n672_), .A2(KEYINPUT111), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n615_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n296_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n722_), .A2(new_n754_), .A3(new_n231_), .A4(new_n652_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT110), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n241_), .A3(new_n515_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g558(.A(G92gat), .B1(new_n752_), .B2(new_n630_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n242_), .A3(new_n629_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n752_), .B2(new_n711_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n594_), .A3(new_n266_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n756_), .A2(new_n254_), .A3(new_n718_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n750_), .A2(new_n718_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n672_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n254_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT113), .B1(new_n672_), .B2(new_n768_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n767_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT53), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n767_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  NAND4_X1  g579(.A1(new_n630_), .A2(new_n515_), .A3(new_n573_), .A4(new_n594_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT118), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n607_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n601_), .B1(new_n596_), .B2(new_n273_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n610_), .B1(new_n605_), .B2(new_n786_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n784_), .A2(new_n610_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n324_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n316_), .B(KEYINPUT55), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n313_), .A2(new_n315_), .A3(new_n314_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n303_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(KEYINPUT115), .A3(new_n303_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n790_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n321_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT117), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n321_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n797_), .B2(KEYINPUT117), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n789_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT58), .B(new_n789_), .C1(new_n798_), .C2(new_n800_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(new_n300_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n611_), .A2(new_n324_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n797_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n799_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n325_), .B2(new_n788_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n325_), .A2(new_n809_), .A3(new_n788_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n296_), .B1(new_n808_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n321_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n611_), .B(new_n324_), .C1(new_n817_), .C2(new_n797_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n325_), .A2(new_n809_), .A3(new_n788_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n810_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT57), .A3(new_n296_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n816_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n231_), .B1(new_n805_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n301_), .A2(new_n673_), .A3(new_n329_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n825_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n783_), .B1(new_n824_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n611_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n296_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n815_), .B(new_n754_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n803_), .A2(new_n300_), .A3(new_n804_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n618_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n830_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n782_), .B(new_n835_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n842_), .B(new_n611_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n833_), .B1(new_n845_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n847_));
  AOI21_X1  g646(.A(G120gat), .B1(new_n652_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n847_), .B2(G120gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n831_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT120), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n842_), .B1(new_n831_), .B2(new_n843_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852_), .B2(new_n329_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n231_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n842_), .B(new_n856_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n618_), .B(new_n782_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n855_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n857_), .A2(KEYINPUT121), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT121), .B1(new_n857_), .B2(new_n859_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  INV_X1    g661(.A(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n831_), .A2(new_n863_), .A3(new_n754_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n842_), .B(new_n300_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n866_), .B2(new_n863_), .ZN(G1343gat));
  NAND3_X1  g666(.A1(new_n630_), .A2(new_n515_), .A3(new_n718_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n711_), .B(new_n869_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n673_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n470_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n329_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n471_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n870_), .A2(new_n231_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n875_), .B(new_n876_), .Z(G1346gat));
  OAI21_X1  g676(.A(new_n462_), .B1(new_n870_), .B2(new_n296_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n824_), .A2(new_n830_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n669_), .A2(new_n462_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n711_), .A3(new_n869_), .A4(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT122), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n878_), .A2(new_n881_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1347gat));
  AOI21_X1  g685(.A(new_n360_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n629_), .A2(new_n573_), .A3(new_n533_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n879_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n889_), .B2(new_n673_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  OAI221_X1 g691(.A(new_n887_), .B1(KEYINPUT123), .B2(KEYINPUT62), .C1(new_n889_), .C2(new_n673_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n889_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n894_), .A2(new_n611_), .A3(new_n449_), .A4(new_n364_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n893_), .A3(new_n895_), .ZN(G1348gat));
  NAND3_X1  g695(.A1(new_n879_), .A2(new_n652_), .A3(new_n888_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(KEYINPUT124), .B2(new_n419_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT124), .B(G176gat), .Z(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(new_n899_), .ZN(G1349gat));
  AND2_X1   g699(.A1(new_n381_), .A2(new_n383_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n373_), .A2(KEYINPUT125), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n894_), .A2(new_n901_), .A3(new_n618_), .A4(new_n902_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n889_), .A2(new_n231_), .B1(KEYINPUT125), .B2(G183gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n889_), .B2(new_n299_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n754_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n889_), .B2(new_n907_), .ZN(G1351gat));
  NAND2_X1  g707(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n630_), .A2(new_n515_), .A3(new_n573_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n711_), .B(new_n910_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n673_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT127), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n912_), .B(new_n914_), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n911_), .A2(new_n329_), .ZN(new_n916_));
  MUX2_X1   g715(.A(G204gat), .B(new_n406_), .S(new_n916_), .Z(G1353gat));
  NOR2_X1   g716(.A1(new_n911_), .A2(new_n231_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n918_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT63), .B(G211gat), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n918_), .B2(new_n920_), .ZN(G1354gat));
  OAI21_X1  g720(.A(G218gat), .B1(new_n911_), .B2(new_n299_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n296_), .A2(G218gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n911_), .B2(new_n923_), .ZN(G1355gat));
endmodule


