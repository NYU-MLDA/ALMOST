//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT95), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT95), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n211_), .B(new_n203_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G183gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT26), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n218_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT79), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G183gat), .A3(G190gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR3_X1    g033(.A1(new_n210_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n213_), .A2(new_n226_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G197gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G204gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n237_), .A2(G204gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT21), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G211gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(G218gat), .ZN(new_n243_));
  INV_X1    g042(.A(G218gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G211gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT87), .B1(new_n237_), .B2(G204gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT87), .ZN(new_n248_));
  INV_X1    g047(.A(G204gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(G197gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n250_), .A3(new_n238_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT88), .B(KEYINPUT21), .Z(new_n252_));
  OAI211_X1 g051(.A(new_n241_), .B(new_n246_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT23), .B1(new_n229_), .B2(new_n231_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n227_), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  OAI22_X1  g054(.A1(new_n254_), .A2(new_n255_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n208_), .A2(KEYINPUT22), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G169gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n257_), .A2(new_n259_), .A3(KEYINPUT96), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT96), .B1(new_n257_), .B2(new_n259_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n209_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(new_n262_), .A3(new_n203_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n244_), .A2(G211gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n242_), .A2(G218gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(KEYINPUT89), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n251_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n247_), .A2(new_n250_), .A3(KEYINPUT90), .A4(new_n238_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n269_), .A2(new_n271_), .A3(KEYINPUT21), .A4(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n236_), .A2(new_n253_), .A3(new_n263_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT97), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n273_), .A2(new_n253_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT97), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n236_), .A4(new_n263_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT19), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n273_), .A2(new_n253_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n232_), .A2(new_n284_), .A3(new_n233_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(new_n208_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n290_), .B2(new_n203_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n216_), .B2(G183gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT26), .B1(new_n219_), .B2(KEYINPUT78), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n221_), .A3(G190gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI22_X1  g099(.A1(new_n285_), .A2(new_n287_), .B1(new_n292_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n282_), .B1(new_n283_), .B2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n275_), .A2(new_n278_), .A3(new_n281_), .A4(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G8gat), .B(G36gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT18), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n301_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n236_), .A2(new_n263_), .B1(new_n253_), .B2(new_n273_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n280_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n303_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n303_), .B2(new_n310_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n202_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT101), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n303_), .A2(new_n310_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n307_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT101), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n202_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT98), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n302_), .A2(new_n274_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n280_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n283_), .A2(new_n301_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n236_), .A2(new_n263_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n283_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT20), .A4(new_n281_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n308_), .A2(new_n309_), .A3(new_n280_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(KEYINPUT98), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n316_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n318_), .A2(KEYINPUT27), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT100), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n281_), .B1(new_n302_), .B2(new_n274_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT98), .B1(new_n331_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(new_n323_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n307_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n318_), .A2(KEYINPUT27), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT100), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n322_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT91), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n283_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G106gat), .ZN(new_n350_));
  INV_X1    g149(.A(G106gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n346_), .A2(new_n351_), .A3(new_n348_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G141gat), .B(G148gat), .Z(new_n353_));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT84), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(G155gat), .A3(G162gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G155gat), .ZN(new_n360_));
  INV_X1    g159(.A(G162gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT83), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT83), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(G155gat), .B2(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n358_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n353_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n369_));
  INV_X1    g168(.A(G141gat), .ZN(new_n370_));
  INV_X1    g169(.A(G148gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n374_));
  OAI22_X1  g173(.A1(KEYINPUT85), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n364_), .A2(new_n362_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n355_), .A2(new_n357_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n365_), .A2(new_n381_), .A3(new_n379_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n368_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT29), .ZN(new_n385_));
  INV_X1    g184(.A(G78gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n283_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n385_), .B2(new_n283_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n350_), .B(new_n352_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n283_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G78gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n351_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n393_));
  AOI211_X1 g192(.A(G106gat), .B(new_n347_), .C1(new_n283_), .C2(new_n345_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n387_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  OR3_X1    g195(.A1(new_n384_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT28), .B1(new_n384_), .B2(KEYINPUT29), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT92), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n398_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n399_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n400_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n396_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n406_), .B2(new_n400_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n413_), .B(KEYINPUT81), .Z(new_n414_));
  AND2_X1   g213(.A1(new_n301_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n301_), .A2(new_n414_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT31), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT31), .B1(new_n415_), .B2(new_n416_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G113gat), .B(G120gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G134gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G127gat), .ZN(new_n430_));
  INV_X1    g229(.A(G127gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G134gat), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT82), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT82), .B1(new_n430_), .B2(new_n432_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n428_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n432_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT82), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n427_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n426_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n421_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n419_), .A2(new_n420_), .A3(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n365_), .A2(new_n381_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT86), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n382_), .A3(new_n377_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n450_), .A2(new_n368_), .B1(new_n440_), .B2(new_n435_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n447_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n384_), .A2(new_n441_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n450_), .A2(new_n440_), .A3(new_n435_), .A4(new_n368_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n455_), .A3(new_n447_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT0), .B(G57gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  AND3_X1   g261(.A1(new_n457_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n412_), .A2(new_n446_), .A3(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n344_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n454_), .A2(new_n455_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n456_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n447_), .B1(new_n454_), .B2(KEYINPUT4), .ZN(new_n474_));
  OAI221_X1 g273(.A(new_n471_), .B1(new_n472_), .B2(new_n447_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n457_), .A2(KEYINPUT33), .A3(new_n458_), .A4(new_n462_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n470_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n307_), .A2(KEYINPUT32), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n303_), .A2(new_n478_), .A3(new_n310_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n477_), .A2(new_n319_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n412_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT99), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n409_), .A2(new_n411_), .A3(new_n465_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n322_), .A2(new_n343_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(KEYINPUT99), .A3(new_n412_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n446_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n467_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  INV_X1    g292(.A(G8gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G1gat), .B(G8gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G43gat), .B(G50gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n498_), .B(new_n501_), .Z(new_n502_));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n501_), .B(KEYINPUT15), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n498_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n498_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n501_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n509_), .A3(new_n503_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G113gat), .B(G141gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n513_), .B(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n491_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT66), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n522_), .A2(KEYINPUT66), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT11), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G71gat), .B(G78gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n522_), .A2(KEYINPUT66), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT11), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n523_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT11), .B(new_n527_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n498_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538_));
  XOR2_X1   g337(.A(G127gat), .B(G155gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G183gat), .B(G211gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n537_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(KEYINPUT17), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(G85gat), .ZN(new_n550_));
  INV_X1    g349(.A(G92gat), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT9), .ZN(new_n552_));
  XOR2_X1   g351(.A(G85gat), .B(G92gat), .Z(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n553_), .B2(KEYINPUT9), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT10), .B(G99gat), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n549_), .B(new_n554_), .C1(G106gat), .C2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n548_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n547_), .A2(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT65), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n547_), .A2(new_n557_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n562_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT65), .B1(new_n565_), .B2(new_n559_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n558_), .A2(new_n563_), .A3(new_n564_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n553_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT8), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n565_), .A2(new_n559_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n568_), .B1(new_n549_), .B2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n556_), .B(new_n571_), .C1(new_n573_), .C2(KEYINPUT8), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n575_), .A2(new_n501_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT68), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n558_), .A2(new_n564_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n572_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n553_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n569_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n586_), .A2(KEYINPUT68), .A3(new_n571_), .A4(new_n556_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n582_), .A2(new_n587_), .A3(new_n506_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n579_), .A2(new_n576_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n580_), .B2(new_n588_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NOR4_X1   g395(.A1(new_n592_), .A2(new_n593_), .A3(KEYINPUT36), .A4(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(KEYINPUT36), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n593_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n600_), .B2(new_n591_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT37), .B1(new_n597_), .B2(new_n601_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n546_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n534_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n574_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n582_), .A2(new_n587_), .A3(KEYINPUT12), .A4(new_n607_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT69), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n612_), .B(new_n613_), .C1(new_n607_), .C2(new_n574_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n534_), .A2(new_n586_), .A3(new_n571_), .A4(new_n556_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n612_), .B1(new_n616_), .B2(new_n613_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n610_), .B(new_n611_), .C1(new_n615_), .C2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n575_), .A2(new_n534_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n613_), .B1(new_n619_), .B2(KEYINPUT67), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT67), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n608_), .A2(new_n616_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(G120gat), .B(G148gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n618_), .A2(new_n623_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT72), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT72), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n618_), .A2(new_n623_), .A3(new_n631_), .A4(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n611_), .A2(new_n610_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n613_), .B1(new_n607_), .B2(new_n574_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT69), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n614_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n634_), .A2(new_n637_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n628_), .B(KEYINPUT71), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n633_), .A2(KEYINPUT13), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT13), .B1(new_n633_), .B2(new_n640_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n521_), .A2(new_n606_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT102), .ZN(new_n646_));
  INV_X1    g445(.A(new_n465_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n493_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT103), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n646_), .A2(new_n650_), .A3(new_n493_), .A4(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT104), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n649_), .A2(new_n655_), .A3(KEYINPUT38), .A4(new_n651_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n491_), .A2(new_n602_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n643_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n641_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n660_), .A2(new_n520_), .A3(new_n546_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n493_), .B1(new_n662_), .B2(new_n647_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n657_), .A2(new_n664_), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n344_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n494_), .B1(KEYINPUT105), .B2(KEYINPUT39), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n668_), .B(new_n669_), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n646_), .A2(new_n494_), .A3(new_n344_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n662_), .B2(new_n446_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT41), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n446_), .A2(new_n674_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n645_), .B2(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n412_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n662_), .B2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT42), .Z(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n679_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n645_), .B2(new_n683_), .ZN(G1327gat));
  AND4_X1   g483(.A1(new_n521_), .A2(new_n602_), .A3(new_n546_), .A4(new_n644_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n647_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n604_), .A2(new_n605_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n491_), .B2(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n491_), .A2(KEYINPUT43), .A3(new_n687_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NOR4_X1   g490(.A1(new_n491_), .A2(KEYINPUT106), .A3(KEYINPUT43), .A4(new_n687_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n546_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n660_), .A2(new_n520_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n695_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n647_), .A2(G29gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n686_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n344_), .A2(KEYINPUT107), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n344_), .A2(KEYINPUT107), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n685_), .A2(new_n703_), .A3(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n708_), .A2(new_n710_), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n711_), .A2(new_n712_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n698_), .A2(new_n344_), .A3(new_n699_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G36gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n715_), .A2(new_n719_), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n718_), .B(new_n713_), .C1(new_n714_), .C2(G36gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  NAND3_X1  g521(.A1(new_n700_), .A2(G43gat), .A3(new_n446_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  AOI21_X1  g523(.A(G43gat), .B1(new_n685_), .B2(new_n446_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n727_));
  AND4_X1   g526(.A1(G43gat), .A2(new_n698_), .A3(new_n446_), .A4(new_n699_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT47), .B1(new_n728_), .B2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  AOI21_X1  g529(.A(G50gat), .B1(new_n685_), .B2(new_n680_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n680_), .A2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n700_), .B2(new_n732_), .ZN(G1331gat));
  NAND4_X1  g532(.A1(new_n658_), .A2(new_n520_), .A3(new_n694_), .A4(new_n660_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n465_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n520_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n491_), .A2(new_n736_), .A3(new_n644_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n606_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n465_), .A2(G57gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1332gat));
  OAI21_X1  g539(.A(G64gat), .B1(new_n734_), .B2(new_n706_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT48), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n706_), .A2(G64gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT110), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n738_), .B2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n734_), .B2(new_n490_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n490_), .A2(G71gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n738_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n734_), .B2(new_n412_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n680_), .A2(new_n386_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n738_), .B2(new_n752_), .ZN(G1335gat));
  NAND3_X1  g552(.A1(new_n660_), .A2(new_n520_), .A3(new_n546_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT112), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n693_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n693_), .A2(KEYINPUT113), .A3(new_n755_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n465_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n737_), .A2(new_n602_), .A3(new_n546_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT111), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n550_), .A3(new_n647_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n760_), .B2(new_n706_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n551_), .A3(new_n344_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1337gat));
  NOR2_X1   g567(.A1(new_n490_), .A2(new_n555_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n763_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n490_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n771_));
  INV_X1    g570(.A(G99gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n770_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n763_), .A2(new_n351_), .A3(new_n680_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n680_), .B(new_n755_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(KEYINPUT52), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(G106gat), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT114), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n787_), .B2(new_n781_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n778_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n778_), .C1(new_n784_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  NAND4_X1  g592(.A1(new_n606_), .A2(new_n659_), .A3(new_n520_), .A4(new_n641_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n795_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n644_), .A2(new_n520_), .A3(new_n606_), .A4(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n796_), .A2(new_n798_), .B1(KEYINPUT115), .B2(KEYINPUT54), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n633_), .A2(new_n640_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n502_), .A2(new_n503_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n507_), .A2(new_n509_), .A3(new_n504_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n519_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n511_), .A2(new_n518_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n618_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n634_), .A2(new_n637_), .A3(KEYINPUT55), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n611_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(G230gat), .A3(G233gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n639_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n813_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n520_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n814_), .A2(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n631_), .B1(new_n638_), .B2(new_n628_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n632_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n736_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(KEYINPUT116), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n806_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n602_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n812_), .A2(new_n813_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n813_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n821_), .A2(KEYINPUT116), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n816_), .A2(new_n817_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n602_), .B1(new_n835_), .B2(new_n806_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n805_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n633_), .B2(new_n805_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n687_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n805_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT117), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n832_), .A2(new_n846_), .A3(KEYINPUT58), .A4(new_n840_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n844_), .A3(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n827_), .A2(new_n837_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n799_), .B1(new_n849_), .B2(new_n546_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n344_), .A2(new_n490_), .A3(new_n465_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n850_), .A2(new_n680_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G113gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n736_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n832_), .A2(new_n846_), .A3(new_n840_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n687_), .B1(new_n857_), .B2(new_n838_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n826_), .A2(new_n825_), .B1(new_n858_), .B2(new_n847_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n694_), .B1(new_n859_), .B2(new_n837_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n412_), .B(new_n851_), .C1(new_n860_), .C2(new_n799_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n856_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n850_), .A2(new_n680_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(KEYINPUT118), .A3(KEYINPUT59), .A4(new_n851_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n520_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n855_), .B1(new_n866_), .B2(new_n854_), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n853_), .B(new_n869_), .C1(KEYINPUT60), .C2(new_n868_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n644_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872_));
  OAI21_X1  g671(.A(G120gat), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT119), .B(new_n644_), .C1(new_n863_), .C2(new_n865_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n870_), .B1(new_n873_), .B2(new_n874_), .ZN(G1341gat));
  OAI21_X1  g674(.A(new_n431_), .B1(new_n861_), .B2(new_n546_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT120), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n431_), .B(new_n546_), .C1(new_n863_), .C2(new_n865_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1342gat));
  NOR2_X1   g678(.A1(new_n687_), .A2(new_n429_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT59), .B1(new_n853_), .B2(KEYINPUT118), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n861_), .A2(new_n862_), .A3(new_n856_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G134gat), .B1(new_n853_), .B2(new_n602_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT121), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n880_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n884_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n886_), .A2(new_n890_), .ZN(G1343gat));
  NOR2_X1   g690(.A1(new_n850_), .A2(new_n446_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n707_), .A2(new_n412_), .A3(new_n465_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n520_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n370_), .ZN(G1344gat));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n644_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n371_), .ZN(G1345gat));
  NOR2_X1   g697(.A1(new_n894_), .A2(new_n546_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT61), .B(G155gat), .Z(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  OAI21_X1  g700(.A(new_n361_), .B1(new_n894_), .B2(new_n824_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n844_), .A2(G162gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT122), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n894_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n902_), .B(KEYINPUT123), .C1(new_n894_), .C2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1347gat));
  OAI21_X1  g708(.A(new_n412_), .B1(new_n860_), .B2(new_n799_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n446_), .A2(new_n465_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n706_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n910_), .A2(new_n913_), .ZN(new_n914_));
  AOI211_X1 g713(.A(KEYINPUT62), .B(new_n208_), .C1(new_n914_), .C2(new_n736_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n736_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(G169gat), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n914_), .B(new_n736_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n915_), .B1(new_n918_), .B2(new_n919_), .ZN(G1348gat));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n864_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n910_), .A2(KEYINPUT124), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n913_), .A2(new_n209_), .A3(new_n644_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G176gat), .B1(new_n914_), .B2(new_n660_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927_));
  OR3_X1    g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1349gat));
  NAND2_X1  g729(.A1(new_n864_), .A2(new_n912_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n931_), .A2(new_n218_), .A3(new_n546_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n922_), .A2(new_n923_), .A3(new_n694_), .A4(new_n912_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n214_), .ZN(G1350gat));
  OAI21_X1  g733(.A(G190gat), .B1(new_n931_), .B2(new_n687_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n224_), .A2(new_n225_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n914_), .A2(new_n936_), .A3(new_n602_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(KEYINPUT126), .ZN(G1351gat));
  NAND3_X1  g738(.A1(new_n892_), .A2(new_n486_), .A3(new_n707_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n520_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n237_), .ZN(G1352gat));
  NOR2_X1   g741(.A1(new_n940_), .A2(new_n644_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n249_), .ZN(G1353gat));
  NOR2_X1   g743(.A1(new_n940_), .A2(new_n546_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n945_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT63), .B(G211gat), .Z(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n945_), .B2(new_n947_), .ZN(G1354gat));
  NOR3_X1   g747(.A1(new_n940_), .A2(new_n244_), .A3(new_n687_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n940_), .A2(new_n824_), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n950_), .A2(KEYINPUT127), .ZN(new_n951_));
  AOI21_X1  g750(.A(G218gat), .B1(new_n950_), .B2(KEYINPUT127), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n949_), .B1(new_n951_), .B2(new_n952_), .ZN(G1355gat));
endmodule


