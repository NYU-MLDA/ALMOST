//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  INV_X1    g000(.A(G134gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G127gat), .ZN(new_n203_));
  INV_X1    g002(.A(G127gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G113gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G120gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(G120gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(new_n203_), .A3(new_n205_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT22), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G169gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n214_), .B1(new_n219_), .B2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT79), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(KEYINPUT79), .B(new_n214_), .C1(new_n219_), .C2(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n222_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n214_), .A2(KEYINPUT24), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  MUX2_X1   g037(.A(new_n237_), .B(KEYINPUT24), .S(new_n238_), .Z(new_n239_));
  AND3_X1   g038(.A1(new_n224_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT78), .B1(new_n224_), .B2(KEYINPUT23), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n227_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT77), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n236_), .A2(new_n239_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n231_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G15gat), .B(G43gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT80), .ZN(new_n247_));
  INV_X1    g046(.A(G71gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(G99gat), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(G99gat), .B1(new_n249_), .B2(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n245_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n231_), .A2(new_n244_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n251_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n213_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT81), .Z(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT30), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT31), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n254_), .A2(new_n257_), .A3(new_n213_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n263_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n258_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G228gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G78gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G106gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G22gat), .B(G50gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G155gat), .ZN(new_n276_));
  INV_X1    g075(.A(G162gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT83), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(G155gat), .B2(G162gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n278_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283_));
  INV_X1    g082(.A(G141gat), .ZN(new_n284_));
  INV_X1    g083(.A(G148gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT2), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n286_), .A2(new_n289_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n282_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n281_), .A2(KEYINPUT1), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(G155gat), .A3(G162gat), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n278_), .A2(new_n294_), .A3(new_n280_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n293_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT28), .B1(new_n304_), .B2(KEYINPUT29), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n292_), .A2(new_n282_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(G197gat), .ZN(new_n313_));
  INV_X1    g112(.A(G197gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT21), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(G197gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n316_), .A2(new_n317_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n314_), .A2(G204gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT84), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI211_X1 g126(.A(KEYINPUT84), .B(new_n317_), .C1(new_n318_), .C2(new_n324_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n322_), .B(new_n323_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n316_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n323_), .A2(new_n317_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n329_), .A2(new_n332_), .B1(new_n304_), .B2(KEYINPUT29), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n310_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n310_), .A2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n275_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n334_), .A3(new_n274_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT33), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n206_), .B(new_n211_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n297_), .A2(new_n302_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n278_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n291_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n290_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n344_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n342_), .B1(new_n343_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n213_), .A2(new_n293_), .A3(new_n303_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT89), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT89), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n306_), .A2(new_n355_), .A3(new_n213_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G57gat), .B(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n306_), .A2(new_n213_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n365_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n359_), .B(new_n364_), .C1(new_n366_), .C2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n341_), .B1(new_n371_), .B2(KEYINPUT91), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT89), .B1(new_n306_), .B2(new_n213_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n213_), .A2(new_n303_), .A3(new_n293_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n356_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT4), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n358_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(KEYINPUT92), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(new_n366_), .B2(new_n378_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n364_), .B1(new_n357_), .B2(new_n369_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n372_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n322_), .A2(new_n323_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n325_), .B(new_n326_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n386_), .A2(new_n387_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n220_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n242_), .A2(KEYINPUT87), .A3(new_n229_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT87), .B1(new_n242_), .B2(new_n229_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n239_), .A2(new_n234_), .A3(new_n228_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT88), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT19), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n329_), .A2(new_n332_), .ZN(new_n399_));
  AOI211_X1 g198(.A(new_n396_), .B(new_n398_), .C1(new_n256_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT88), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n388_), .A2(new_n392_), .A3(new_n401_), .A4(new_n393_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n392_), .A2(new_n393_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n256_), .B2(new_n399_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n398_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n403_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n407_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n371_), .A2(KEYINPUT91), .A3(new_n341_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n385_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n403_), .A2(new_n410_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n407_), .A2(KEYINPUT32), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n359_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n364_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n371_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n396_), .B1(new_n256_), .B2(new_n399_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n394_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n398_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n392_), .A2(new_n393_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n399_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n396_), .B1(new_n245_), .B2(new_n388_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n398_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n417_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n423_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AOI211_X1 g233(.A(KEYINPUT93), .B(new_n417_), .C1(new_n426_), .C2(new_n431_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n418_), .B(new_n422_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n340_), .B1(new_n415_), .B2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n403_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n407_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n408_), .A2(new_n409_), .A3(new_n398_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n430_), .B1(new_n394_), .B2(new_n424_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n442_), .A3(KEYINPUT27), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT94), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT94), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n438_), .A2(new_n442_), .A3(new_n447_), .A4(KEYINPUT27), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n340_), .A2(new_n421_), .A3(new_n371_), .ZN(new_n449_));
  AND4_X1   g248(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n269_), .B1(new_n437_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT95), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n446_), .A2(new_n448_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n454_), .A2(new_n444_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n340_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n269_), .A2(new_n422_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(KEYINPUT95), .B(new_n269_), .C1(new_n437_), .C2(new_n450_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT68), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n463_), .A2(KEYINPUT68), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(KEYINPUT68), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT71), .B(G1gat), .ZN(new_n473_));
  INV_X1    g272(.A(G8gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT14), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n475_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n471_), .B1(new_n481_), .B2(new_n480_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n462_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT74), .ZN(new_n486_));
  INV_X1    g285(.A(new_n484_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n461_), .B(new_n487_), .C1(new_n488_), .C2(new_n482_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n490_), .B(new_n462_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n493_));
  XOR2_X1   g292(.A(G113gat), .B(G141gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT75), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G169gat), .B(G197gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n460_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G85gat), .B(G92gat), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT9), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT10), .B(G99gat), .ZN(new_n507_));
  OAI221_X1 g306(.A(new_n505_), .B1(KEYINPUT9), .B2(new_n506_), .C1(G106gat), .C2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT7), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n504_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n516_), .B2(new_n504_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n513_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT34), .ZN(new_n522_));
  OAI22_X1  g321(.A1(new_n520_), .A2(new_n471_), .B1(KEYINPUT35), .B2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n508_), .A2(new_n512_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n516_), .A2(new_n504_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT8), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n516_), .A2(new_n517_), .A3(new_n504_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n488_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n522_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n523_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n532_), .B1(new_n523_), .B2(new_n529_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n536_), .B(KEYINPUT36), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT70), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n543_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(new_n545_), .A3(new_n539_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n539_), .A2(KEYINPUT69), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n533_), .A2(new_n552_), .A3(new_n537_), .A4(new_n538_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n546_), .A2(new_n550_), .B1(KEYINPUT37), .B2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT65), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n560_));
  XOR2_X1   g359(.A(G71gat), .B(G78gat), .Z(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n560_), .A2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n557_), .B1(new_n520_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n528_), .A2(KEYINPUT65), .A3(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n528_), .A2(new_n564_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n556_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n571_));
  NOR2_X1   g370(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n572_));
  OAI22_X1  g371(.A1(new_n528_), .A2(new_n564_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n520_), .B(new_n565_), .C1(KEYINPUT66), .C2(KEYINPUT12), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n556_), .B1(new_n528_), .B2(new_n564_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G120gat), .B(G148gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n570_), .A2(new_n576_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(KEYINPUT13), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT17), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(KEYINPUT72), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n564_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n482_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(KEYINPUT73), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n602_), .B2(new_n594_), .ZN(new_n603_));
  AOI211_X1 g402(.A(new_n595_), .B(new_n597_), .C1(new_n600_), .C2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n601_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n555_), .A2(new_n590_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n503_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(new_n422_), .A3(new_n473_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n544_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n460_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n590_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n502_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n608_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n422_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n612_), .A2(new_n613_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n614_), .A2(new_n622_), .A3(new_n623_), .ZN(G1324gat));
  OAI21_X1  g423(.A(G8gat), .B1(new_n620_), .B2(new_n455_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n454_), .A2(new_n444_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n611_), .A2(new_n474_), .A3(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g429(.A(G15gat), .B1(new_n620_), .B2(new_n269_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT96), .B(KEYINPUT41), .Z(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n610_), .A2(G15gat), .A3(new_n269_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n633_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n620_), .B2(new_n456_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n456_), .A2(G22gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n610_), .B2(new_n640_), .ZN(G1327gat));
  NAND2_X1  g440(.A1(new_n544_), .A2(new_n608_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n590_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n503_), .A2(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n644_), .A2(G29gat), .A3(new_n621_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n618_), .A2(new_n607_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n458_), .A2(new_n459_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n371_), .A2(KEYINPUT91), .A3(new_n341_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n650_), .A2(new_n372_), .A3(new_n384_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n433_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT93), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n432_), .A2(new_n423_), .A3(new_n433_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n416_), .A2(new_n417_), .B1(new_n421_), .B2(new_n371_), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n651_), .A2(new_n413_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n649_), .B1(new_n657_), .B2(new_n340_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT95), .B1(new_n658_), .B2(new_n269_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n647_), .B(new_n555_), .C1(new_n648_), .C2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT97), .B(KEYINPUT43), .Z(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n460_), .B2(new_n555_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n646_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n646_), .C1(new_n661_), .C2(new_n664_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n422_), .A3(new_n668_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(KEYINPUT98), .A3(G29gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT98), .B1(new_n669_), .B2(G29gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n645_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  NAND2_X1  g471(.A1(new_n455_), .A2(KEYINPUT100), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n627_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n644_), .A2(G36gat), .A3(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT45), .Z(new_n679_));
  NAND3_X1  g478(.A1(new_n667_), .A2(new_n627_), .A3(new_n668_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT99), .A3(G36gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT99), .B1(new_n680_), .B2(G36gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n679_), .B(KEYINPUT46), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  INV_X1    g486(.A(new_n269_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n667_), .A2(G43gat), .A3(new_n688_), .A4(new_n668_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n644_), .A2(new_n269_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(G43gat), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g491(.A1(new_n644_), .A2(G50gat), .A3(new_n456_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n667_), .A2(new_n340_), .A3(new_n668_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(KEYINPUT101), .A3(G50gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT101), .B1(new_n694_), .B2(G50gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1331gat));
  NAND4_X1  g496(.A1(new_n616_), .A2(new_n501_), .A3(new_n590_), .A4(new_n607_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n621_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n460_), .A2(new_n501_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n546_), .A2(new_n550_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n608_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n590_), .A3(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT102), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n621_), .A2(G57gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n699_), .B1(new_n705_), .B2(new_n706_), .ZN(G1332gat));
  OAI21_X1  g506(.A(G64gat), .B1(new_n698_), .B2(new_n677_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT48), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n677_), .A2(G64gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n705_), .B2(new_n710_), .ZN(G1333gat));
  OAI21_X1  g510(.A(G71gat), .B1(new_n698_), .B2(new_n269_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT49), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n688_), .A2(new_n248_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n705_), .B2(new_n714_), .ZN(G1334gat));
  OAI21_X1  g514(.A(G78gat), .B1(new_n698_), .B2(new_n456_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT103), .Z(new_n717_));
  OR2_X1    g516(.A1(new_n717_), .A2(KEYINPUT50), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(KEYINPUT50), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n705_), .A2(G78gat), .A3(new_n456_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n720_), .ZN(G1335gat));
  NAND2_X1  g520(.A1(new_n460_), .A2(new_n555_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n662_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n660_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(KEYINPUT104), .A3(new_n660_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n590_), .A2(new_n501_), .A3(new_n608_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n727_), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730_), .B2(new_n621_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n700_), .A2(new_n590_), .A3(new_n608_), .A4(new_n544_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n621_), .A2(G85gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n732_), .B2(new_n733_), .ZN(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n730_), .B2(new_n677_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n455_), .A2(G92gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n732_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1337gat));
  AND2_X1   g538(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n732_), .A2(new_n269_), .A3(new_n507_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n726_), .A2(new_n688_), .A3(new_n727_), .A4(new_n729_), .ZN(new_n742_));
  AOI211_X1 g541(.A(new_n740_), .B(new_n741_), .C1(new_n742_), .C2(G99gat), .ZN(new_n743_));
  NOR2_X1   g542(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1338gat));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n456_), .B(new_n728_), .C1(new_n723_), .C2(new_n660_), .ZN(new_n747_));
  INV_X1    g546(.A(G106gat), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n747_), .A2(KEYINPUT108), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n724_), .A2(new_n340_), .A3(new_n729_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G106gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n746_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n732_), .A2(G106gat), .A3(new_n456_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT107), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT108), .B1(new_n747_), .B2(new_n748_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n751_), .A2(new_n750_), .A3(G106gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(KEYINPUT52), .A3(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n753_), .A2(new_n755_), .A3(new_n761_), .A4(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  NAND2_X1  g562(.A1(new_n455_), .A2(new_n456_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n688_), .A2(new_n422_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n767_));
  INV_X1    g566(.A(new_n577_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n497_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n486_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(KEYINPUT76), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n768_), .A2(new_n584_), .B1(new_n771_), .B2(new_n498_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n573_), .A2(new_n574_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n556_), .B1(new_n773_), .B2(new_n568_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n576_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .A4(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n582_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n582_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n772_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT110), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n772_), .B(new_n783_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n487_), .B1(new_n488_), .B2(new_n482_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n461_), .B1(new_n785_), .B2(KEYINPUT111), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(KEYINPUT111), .B2(new_n785_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n483_), .A2(new_n484_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n769_), .B1(new_n788_), .B2(new_n461_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(KEYINPUT112), .A3(new_n789_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n792_), .A2(new_n793_), .B1(new_n770_), .B2(new_n769_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n586_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n782_), .A2(new_n784_), .A3(new_n795_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n796_), .A2(KEYINPUT57), .A3(new_n615_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n796_), .B2(new_n615_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n582_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT113), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n778_), .A2(new_n802_), .A3(KEYINPUT56), .A4(new_n582_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n778_), .A2(new_n582_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n585_), .A3(new_n794_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n585_), .A4(new_n794_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n555_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n607_), .B1(new_n799_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT70), .B1(new_n544_), .B2(new_n545_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n548_), .A2(new_n549_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n702_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(new_n501_), .A3(new_n617_), .A4(new_n607_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n703_), .A2(new_n501_), .A3(new_n617_), .A4(new_n818_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n766_), .B(new_n767_), .C1(new_n813_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n766_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n585_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n806_), .B2(new_n800_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n795_), .B1(new_n826_), .B2(new_n783_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n784_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n615_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n796_), .A2(KEYINPUT57), .A3(new_n615_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n812_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n831_), .A2(KEYINPUT114), .A3(new_n812_), .A4(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n608_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n822_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n824_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n823_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n501_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n207_), .A3(new_n502_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1340gat));
  OAI211_X1 g643(.A(new_n590_), .B(new_n823_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(G120gat), .ZN(new_n846_));
  INV_X1    g645(.A(new_n839_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G120gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n617_), .A2(KEYINPUT60), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n847_), .B2(new_n851_), .ZN(G1341gat));
  OAI21_X1  g651(.A(G127gat), .B1(new_n841_), .B2(new_n608_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n822_), .A2(new_n204_), .A3(new_n607_), .A4(new_n766_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1342gat));
  OAI21_X1  g654(.A(G134gat), .B1(new_n841_), .B2(new_n816_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n839_), .A2(new_n202_), .A3(new_n544_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1343gat));
  AOI21_X1  g657(.A(new_n688_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n676_), .A2(new_n456_), .A3(new_n621_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n502_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n590_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n607_), .A3(new_n860_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  AND4_X1   g666(.A1(G162gat), .A2(new_n859_), .A3(new_n555_), .A4(new_n860_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT114), .B1(new_n799_), .B2(new_n812_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n836_), .A2(new_n608_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n838_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(new_n269_), .A3(new_n544_), .A4(new_n860_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n277_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT116), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n875_), .A3(new_n277_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n868_), .B1(new_n874_), .B2(new_n876_), .ZN(G1347gat));
  AND2_X1   g676(.A1(new_n676_), .A2(new_n457_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n502_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT117), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n456_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n822_), .B1(new_n833_), .B2(new_n608_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G169gat), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT62), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n878_), .A2(new_n456_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n885_), .B(new_n887_), .C1(new_n813_), .C2(new_n822_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT118), .B1(new_n882_), .B2(new_n886_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n501_), .A2(new_n219_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT119), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n884_), .A2(new_n893_), .ZN(G1348gat));
  AND4_X1   g693(.A1(G176gat), .A2(new_n871_), .A3(new_n590_), .A4(new_n887_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n888_), .A2(new_n889_), .A3(new_n590_), .ZN(new_n896_));
  INV_X1    g695(.A(G176gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT120), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n900_), .A3(new_n897_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n895_), .B1(new_n899_), .B2(new_n901_), .ZN(G1349gat));
  NOR2_X1   g701(.A1(new_n608_), .A2(new_n232_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n888_), .A2(new_n889_), .A3(new_n903_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n838_), .A2(new_n608_), .A3(new_n886_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n905_), .A2(G183gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT121), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n909_), .A3(new_n906_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1350gat));
  NAND2_X1  g710(.A1(new_n544_), .A2(new_n233_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT123), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n890_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n888_), .A2(new_n889_), .A3(new_n555_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n915_), .A2(new_n916_), .A3(G190gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n915_), .B2(G190gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n914_), .B1(new_n917_), .B2(new_n918_), .ZN(G1351gat));
  NAND2_X1  g718(.A1(new_n676_), .A2(new_n449_), .ZN(new_n920_));
  AOI211_X1 g719(.A(new_n688_), .B(new_n920_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(G197gat), .A4(new_n502_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n920_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n871_), .A2(new_n269_), .A3(new_n502_), .A4(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT124), .B1(new_n925_), .B2(new_n314_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n314_), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n923_), .A2(new_n926_), .A3(new_n927_), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n921_), .A2(new_n590_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(G204gat), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n921_), .B(new_n590_), .C1(KEYINPUT125), .C2(new_n312_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1353gat));
  AOI21_X1  g732(.A(new_n608_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n871_), .A2(new_n269_), .A3(new_n924_), .A4(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n936_), .A2(KEYINPUT126), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n936_), .B(KEYINPUT126), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n935_), .B2(new_n939_), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n921_), .A2(new_n941_), .A3(new_n544_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n921_), .A2(new_n555_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n941_), .ZN(G1355gat));
endmodule


