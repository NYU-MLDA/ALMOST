//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(G57gat), .B(G64gat), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G57gat), .B(G64gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n204_), .A3(KEYINPUT11), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n218_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n213_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n233_), .A2(new_n236_), .A3(new_n223_), .A4(new_n219_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n218_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n216_), .A2(new_n228_), .A3(new_n217_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n237_), .B2(KEYINPUT64), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n222_), .A2(new_n243_), .A3(new_n226_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n229_), .A2(new_n240_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT10), .B(G99gat), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n232_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n247_), .A2(new_n249_), .A3(new_n250_), .A4(new_n226_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n212_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n251_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n257_), .A2(new_n213_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n258_), .B2(new_n240_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT67), .B(new_n255_), .C1(new_n259_), .C2(new_n212_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(KEYINPUT12), .ZN(new_n261_));
  AND2_X1   g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n259_), .B2(new_n212_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n254_), .A2(new_n260_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n212_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n266_), .B2(new_n252_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT69), .ZN(new_n270_));
  XOR2_X1   g069(.A(G120gat), .B(G148gat), .Z(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n268_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n264_), .A2(new_n267_), .A3(new_n274_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n268_), .A2(KEYINPUT70), .A3(new_n275_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n284_), .A2(KEYINPUT71), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n282_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n288_), .B(new_n289_), .C1(new_n281_), .C2(new_n285_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G50gat), .ZN(new_n299_));
  INV_X1    g098(.A(G36gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G29gat), .ZN(new_n301_));
  INV_X1    g100(.A(G29gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G36gat), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n301_), .A2(new_n303_), .A3(KEYINPUT75), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT75), .B1(new_n301_), .B2(new_n303_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n304_), .A2(new_n305_), .A3(G43gat), .ZN(new_n306_));
  INV_X1    g105(.A(G43gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n302_), .A2(G36gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n300_), .A2(G29gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n301_), .A2(new_n303_), .A3(KEYINPUT75), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n307_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n299_), .B1(new_n306_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(G43gat), .B1(new_n304_), .B2(new_n305_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(G50gat), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n314_), .A2(KEYINPUT15), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT15), .B1(new_n314_), .B2(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n298_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G229gat), .A2(G233gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT82), .Z(new_n322_));
  AND3_X1   g121(.A1(new_n315_), .A2(G50gat), .A3(new_n316_), .ZN(new_n323_));
  AOI21_X1  g122(.A(G50gat), .B1(new_n315_), .B2(new_n316_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n297_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n296_), .B(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n298_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n314_), .A2(new_n327_), .A3(new_n317_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n321_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT81), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335_));
  AOI211_X1 g134(.A(new_n335_), .B(new_n321_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n329_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G169gat), .B(G197gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT83), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G141gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n329_), .B(new_n341_), .C1(new_n334_), .C2(new_n336_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(KEYINPUT84), .A3(new_n342_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n292_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT23), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  INV_X1    g155(.A(G176gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT25), .B(G183gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT24), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(G169gat), .B2(G176gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n360_), .A2(new_n361_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n362_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n351_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G204gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(G197gat), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(G204gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT21), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n369_), .B2(G197gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n376_), .B(new_n377_), .C1(new_n371_), .C2(G204gat), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n373_), .B(new_n374_), .C1(new_n378_), .C2(KEYINPUT21), .ZN(new_n379_));
  INV_X1    g178(.A(new_n374_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(KEYINPUT21), .A3(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n359_), .A2(new_n368_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n356_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n356_), .A2(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n357_), .A3(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n351_), .A2(new_n353_), .B1(G169gat), .B2(G176gat), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n351_), .A2(new_n367_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n386_), .A2(new_n387_), .B1(new_n388_), .B2(new_n366_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n379_), .A2(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT20), .B(new_n382_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT19), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(KEYINPUT20), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n359_), .A2(new_n368_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(new_n390_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n392_), .A2(new_n395_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT18), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G64gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(new_n215_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT27), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n390_), .A2(KEYINPUT92), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n379_), .A2(new_n408_), .A3(new_n381_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n389_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT20), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT99), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n398_), .A2(new_n390_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n414_), .A3(KEYINPUT20), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n395_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n392_), .A2(new_n395_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n403_), .B(G92gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n392_), .A2(new_n395_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n396_), .A2(new_n399_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n404_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n426_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n429_), .A2(new_n423_), .A3(new_n421_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n428_), .A2(KEYINPUT27), .A3(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n422_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT89), .ZN(new_n435_));
  INV_X1    g234(.A(G155gat), .ZN(new_n436_));
  INV_X1    g235(.A(G162gat), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n435_), .A2(KEYINPUT1), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT90), .B1(new_n435_), .B2(KEYINPUT1), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT89), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n434_), .B(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n438_), .A2(new_n439_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G141gat), .A2(G148gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT88), .ZN(new_n447_));
  INV_X1    g246(.A(G141gat), .ZN(new_n448_));
  INV_X1    g247(.A(G148gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G127gat), .B(G134gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G120gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n448_), .A2(new_n449_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n455_), .A2(KEYINPUT2), .B1(new_n456_), .B2(KEYINPUT3), .ZN(new_n457_));
  OAI221_X1 g256(.A(new_n457_), .B1(KEYINPUT3), .B2(new_n456_), .C1(new_n447_), .C2(KEYINPUT2), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n441_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n454_), .B(KEYINPUT86), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n445_), .A2(new_n450_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n461_), .B(KEYINPUT4), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n462_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n451_), .A2(new_n460_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n433_), .B1(new_n464_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G29gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G85gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n433_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n465_), .A2(new_n466_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(new_n461_), .ZN(new_n478_));
  OR3_X1    g277(.A1(new_n469_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n469_), .B2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n463_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G22gat), .B(G50gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT28), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G78gat), .B(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n407_), .A2(new_n409_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n483_), .B2(new_n463_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n466_), .A2(KEYINPUT29), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n391_), .A2(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n489_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT93), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n487_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n492_), .B1(new_n495_), .B2(new_n490_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n488_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n491_), .A2(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n489_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(new_n505_), .A3(new_n499_), .A4(new_n487_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G15gat), .B(G43gat), .Z(new_n509_));
  XOR2_X1   g308(.A(new_n462_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT30), .B1(new_n359_), .B2(new_n368_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n359_), .A2(new_n368_), .A3(KEYINPUT30), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n514_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n517_), .B1(new_n520_), .B2(new_n512_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n511_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n526_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(new_n510_), .A3(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n507_), .A2(new_n508_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n432_), .B(new_n482_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(KEYINPUT33), .B(new_n475_), .C1(new_n469_), .C2(new_n478_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n477_), .A2(new_n476_), .A3(new_n461_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n535_), .A2(new_n474_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n464_), .A2(new_n433_), .A3(new_n468_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n534_), .B(new_n538_), .C1(new_n428_), .C2(new_n430_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT98), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n480_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n480_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n420_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n429_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n543_), .A2(new_n544_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n508_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT93), .B1(new_n504_), .B2(new_n489_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n551_), .A2(new_n487_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n530_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n533_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n212_), .B(new_n327_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n559_), .A2(KEYINPUT17), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(KEYINPUT79), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n565_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT80), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n556_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n246_), .A2(new_n251_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n259_), .A2(new_n325_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT73), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT35), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(KEYINPUT35), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT74), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n582_), .A2(new_n574_), .A3(new_n575_), .A4(new_n579_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n586_), .A3(new_n590_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT100), .Z(new_n599_));
  NOR2_X1   g398(.A1(new_n572_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n349_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n202_), .B1(new_n601_), .B2(new_n481_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT101), .Z(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n594_), .A2(new_n593_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n587_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n605_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n596_), .A2(new_n597_), .A3(new_n604_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n348_), .B(KEYINPUT85), .Z(new_n612_));
  NOR4_X1   g411(.A1(new_n292_), .A2(new_n572_), .A3(new_n611_), .A4(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n202_), .A3(new_n481_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT38), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n603_), .A2(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n429_), .A2(new_n421_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n423_), .A3(new_n405_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n424_), .A2(new_n427_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT27), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n404_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n623_), .B2(new_n406_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n601_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT102), .B1(new_n625_), .B2(G8gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n630_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n432_), .A2(G8gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n613_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n617_), .B1(new_n631_), .B2(new_n635_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n629_), .A2(new_n630_), .B1(new_n613_), .B2(new_n633_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n629_), .A2(new_n630_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT40), .B(new_n637_), .C1(new_n638_), .C2(new_n628_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(G1325gat));
  INV_X1    g439(.A(G15gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n530_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n601_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n613_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n601_), .B2(new_n553_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT42), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n613_), .A2(new_n647_), .A3(new_n553_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n480_), .A2(new_n541_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT98), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n619_), .A2(new_n620_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n544_), .A4(new_n534_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n548_), .A2(new_n546_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n553_), .A2(new_n642_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n642_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n507_), .A2(new_n508_), .A3(new_n530_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n624_), .A2(new_n481_), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n657_), .A2(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n598_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n663_), .A2(new_n571_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n612_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(new_n291_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n302_), .A3(new_n481_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n663_), .B2(new_n610_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n556_), .A2(KEYINPUT43), .A3(new_n611_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n571_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n292_), .A3(new_n348_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT44), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT103), .B1(new_n677_), .B2(new_n482_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G29gat), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n677_), .A2(KEYINPUT103), .A3(new_n482_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n668_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  OAI21_X1  g480(.A(G36gat), .B1(new_n677_), .B2(new_n432_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n300_), .A3(new_n624_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1329gat));
  NOR3_X1   g486(.A1(new_n677_), .A2(new_n307_), .A3(new_n530_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n667_), .A2(new_n642_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT105), .A3(new_n307_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n689_), .B2(new_n307_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n688_), .A2(KEYINPUT47), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT47), .B1(new_n688_), .B2(new_n692_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1330gat));
  NOR3_X1   g494(.A1(new_n677_), .A2(new_n299_), .A3(new_n554_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G50gat), .B1(new_n667_), .B2(new_n553_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1331gat));
  NAND3_X1  g497(.A1(new_n600_), .A2(new_n292_), .A3(new_n612_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G57gat), .B1(new_n699_), .B2(new_n482_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n287_), .A2(new_n290_), .A3(new_n348_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n701_), .A2(new_n572_), .A3(new_n611_), .ZN(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n481_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n704_), .ZN(G1332gat));
  OAI21_X1  g504(.A(G64gat), .B1(new_n699_), .B2(new_n432_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT48), .ZN(new_n707_));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n708_), .A3(new_n624_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(G1333gat));
  OAI21_X1  g509(.A(G71gat), .B1(new_n699_), .B2(new_n530_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT49), .ZN(new_n712_));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n702_), .A2(new_n713_), .A3(new_n642_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT106), .ZN(G1334gat));
  OAI21_X1  g515(.A(G78gat), .B1(new_n699_), .B2(new_n554_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT50), .ZN(new_n718_));
  INV_X1    g517(.A(G78gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n702_), .A2(new_n719_), .A3(new_n553_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT107), .Z(G1335gat));
  AND3_X1   g521(.A1(new_n287_), .A2(new_n290_), .A3(new_n348_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n665_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n214_), .A3(new_n481_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT108), .B1(new_n673_), .B2(new_n701_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n556_), .A2(new_n611_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n571_), .B1(new_n727_), .B2(new_n669_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(new_n723_), .A3(new_n729_), .A4(new_n671_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n482_), .B1(new_n726_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n731_), .B2(new_n214_), .ZN(G1336gat));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n215_), .A3(new_n624_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n432_), .B1(new_n726_), .B2(new_n730_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n215_), .ZN(G1337gat));
  NAND3_X1  g534(.A1(new_n724_), .A2(new_n248_), .A3(new_n642_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n530_), .B1(new_n726_), .B2(new_n730_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n231_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT109), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(new_n736_), .C1(new_n737_), .C2(new_n231_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(KEYINPUT51), .A3(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n743_));
  OR2_X1    g542(.A1(new_n738_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT111), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1338gat));
  NAND3_X1  g548(.A1(new_n724_), .A2(new_n232_), .A3(new_n553_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n728_), .A2(new_n723_), .A3(new_n553_), .A4(new_n671_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(G106gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G106gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  INV_X1    g556(.A(new_n278_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n320_), .A2(new_n331_), .A3(new_n322_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n322_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n341_), .B1(new_n332_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n345_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n757_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n763_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT115), .A3(new_n278_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n255_), .B1(new_n259_), .B2(new_n212_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n768_), .A2(new_n203_), .B1(KEYINPUT12), .B2(new_n252_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT55), .A3(new_n260_), .A4(new_n263_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n254_), .A2(new_n265_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n262_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n264_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n275_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n767_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n767_), .B(KEYINPUT58), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n611_), .A3(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n279_), .A2(new_n280_), .A3(new_n765_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n775_), .A2(new_n275_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(KEYINPUT113), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n346_), .A2(new_n278_), .A3(new_n347_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n346_), .A2(KEYINPUT112), .A3(new_n278_), .A4(new_n347_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n786_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n784_), .A2(new_n785_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n783_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n664_), .A2(KEYINPUT57), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n782_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n783_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n786_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n776_), .A2(new_n777_), .A3(KEYINPUT113), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n800_), .B1(new_n804_), .B2(new_n664_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(new_n798_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n797_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n610_), .B1(new_n779_), .B2(new_n778_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n804_), .A2(new_n807_), .B1(new_n808_), .B2(new_n781_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n799_), .B1(new_n796_), .B2(new_n598_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n812_), .A3(new_n672_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n288_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(new_n571_), .A3(new_n610_), .A4(new_n612_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n432_), .A2(new_n481_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n659_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n348_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n571_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n817_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n826_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n821_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n831_), .B2(new_n822_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n666_), .A2(G113gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT118), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n824_), .B1(new_n836_), .B2(new_n838_), .ZN(G1340gat));
  OAI21_X1  g638(.A(G120gat), .B1(new_n835_), .B2(new_n291_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n291_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n822_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n835_), .B2(new_n672_), .ZN(new_n845_));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n822_), .A2(new_n846_), .A3(new_n571_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n822_), .B2(new_n599_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n611_), .A2(G134gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT119), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n836_), .B2(new_n851_), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n820_), .A2(new_n660_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n819_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n348_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n448_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n291_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT120), .B(G148gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1345gat));
  NOR2_X1   g658(.A1(new_n854_), .A2(new_n672_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT121), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n860_), .B(new_n862_), .ZN(G1346gat));
  OAI21_X1  g662(.A(G162gat), .B1(new_n854_), .B2(new_n610_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n599_), .A2(new_n437_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n854_), .B2(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g666(.A1(new_n432_), .A2(new_n481_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n659_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n823_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G169gat), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n384_), .A2(new_n385_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n876_), .B(new_n877_), .C1(new_n878_), .C2(new_n873_), .ZN(G1348gat));
  AOI21_X1  g678(.A(G176gat), .B1(new_n872_), .B2(new_n292_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n804_), .A2(new_n807_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n795_), .A2(new_n786_), .A3(new_n789_), .A4(new_n790_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n598_), .B1(new_n882_), .B2(new_n801_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n881_), .B(new_n782_), .C1(new_n883_), .C2(new_n800_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n571_), .B1(new_n884_), .B2(KEYINPUT116), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n817_), .B1(new_n885_), .B2(new_n812_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n553_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n291_), .A2(new_n357_), .A3(new_n530_), .A4(new_n869_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n880_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NAND4_X1  g688(.A1(new_n887_), .A2(new_n571_), .A3(new_n642_), .A4(new_n868_), .ZN(new_n890_));
  INV_X1    g689(.A(G183gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n672_), .A2(new_n360_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n890_), .A2(new_n891_), .B1(new_n872_), .B2(new_n892_), .ZN(G1350gat));
  INV_X1    g692(.A(new_n872_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G190gat), .B1(new_n894_), .B2(new_n610_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n599_), .A2(new_n361_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT123), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n894_), .B2(new_n897_), .ZN(G1351gat));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n869_), .A2(new_n660_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n886_), .B2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n819_), .A2(KEYINPUT124), .A3(new_n900_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n823_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n291_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n369_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT124), .B1(new_n819_), .B2(new_n900_), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n899_), .B(new_n901_), .C1(new_n813_), .C2(new_n818_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n292_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(KEYINPUT125), .A3(G204gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n369_), .B(new_n292_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n904_), .A2(KEYINPUT126), .A3(new_n369_), .A4(new_n292_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n914_), .A2(new_n919_), .ZN(G1353gat));
  NAND2_X1  g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n904_), .A2(new_n571_), .A3(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT127), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n922_), .B(new_n925_), .ZN(G1354gat));
  INV_X1    g725(.A(new_n904_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G218gat), .B1(new_n927_), .B2(new_n610_), .ZN(new_n928_));
  INV_X1    g727(.A(G218gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n904_), .A2(new_n929_), .A3(new_n599_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1355gat));
endmodule


