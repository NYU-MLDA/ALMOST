//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G231gat), .A2(G233gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G71gat), .B(G78gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT11), .ZN(new_n215_));
  INV_X1    g014(.A(new_n214_), .ZN(new_n216_));
  INV_X1    g015(.A(G64gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(G57gat), .ZN(new_n218_));
  INV_X1    g017(.A(G57gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G64gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n220_), .A3(KEYINPUT11), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n215_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n212_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G127gat), .B(G155gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT16), .ZN(new_n228_));
  XOR2_X1   g027(.A(G183gat), .B(G211gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n225_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n225_), .B(KEYINPUT70), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(KEYINPUT17), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT71), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT71), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n231_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G29gat), .B(G36gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT15), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n246_), .A3(new_n210_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n210_), .A2(new_n243_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n248_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT72), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n257_), .A2(KEYINPUT73), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G169gat), .B(G197gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(KEYINPUT73), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n259_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n255_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n250_), .B(new_n254_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT6), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(G99gat), .A3(G106gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n274_));
  INV_X1    g073(.A(G106gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G85gat), .ZN(new_n278_));
  INV_X1    g077(.A(G92gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(KEYINPUT9), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT9), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n273_), .A2(new_n277_), .A3(new_n282_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n281_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI211_X1 g090(.A(KEYINPUT8), .B(new_n287_), .C1(new_n291_), .C2(new_n273_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT8), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n294_));
  INV_X1    g093(.A(G99gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n275_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n273_), .A2(new_n288_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n286_), .B(new_n224_), .C1(new_n292_), .C2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT64), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n270_), .A2(new_n272_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n288_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n298_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT8), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n297_), .A2(new_n293_), .A3(new_n298_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n308_), .A2(KEYINPUT64), .A3(new_n286_), .A4(new_n224_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n286_), .B1(new_n292_), .B2(new_n299_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n224_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G230gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT12), .ZN(new_n318_));
  INV_X1    g117(.A(new_n286_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n320_), .B2(new_n224_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n316_), .B1(new_n320_), .B2(new_n224_), .ZN(new_n322_));
  OAI211_X1 g121(.A(KEYINPUT12), .B(new_n215_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n292_), .A2(new_n299_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n286_), .A2(KEYINPUT65), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n270_), .A2(new_n272_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n277_), .A4(new_n282_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n324_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n322_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n326_), .B(new_n329_), .C1(new_n292_), .C2(new_n299_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n313_), .A2(new_n318_), .B1(new_n335_), .B2(new_n324_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT66), .A3(new_n322_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n317_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G120gat), .B(G148gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT5), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n340_), .B(new_n341_), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n342_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n317_), .A2(new_n334_), .A3(new_n337_), .A4(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n343_), .A2(KEYINPUT13), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT13), .B1(new_n343_), .B2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n237_), .A2(new_n268_), .A3(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT96), .Z(new_n350_));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT91), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n354_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  OR2_X1    g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n359_), .A2(KEYINPUT3), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OR3_X1    g164(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n364_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n362_), .A2(new_n365_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(KEYINPUT1), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT78), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n369_), .A2(KEYINPUT1), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n369_), .A2(new_n376_), .A3(KEYINPUT1), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .A4(new_n371_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G127gat), .B(G134gat), .Z(new_n381_));
  XOR2_X1   g180(.A(G113gat), .B(G120gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(KEYINPUT89), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n372_), .A2(new_n383_), .A3(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT4), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n380_), .A2(KEYINPUT89), .A3(new_n388_), .A4(new_n384_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n358_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n358_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n384_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(new_n386_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n357_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n394_), .A2(KEYINPUT92), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT92), .B1(new_n394_), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(G8gat), .B(G36gat), .Z(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT85), .B(G204gat), .ZN(new_n405_));
  INV_X1    g204(.A(G197gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT83), .B(G197gat), .ZN(new_n408_));
  INV_X1    g207(.A(G204gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT86), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412_));
  OAI221_X1 g211(.A(new_n412_), .B1(new_n408_), .B2(new_n409_), .C1(new_n406_), .C2(new_n405_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G211gat), .B(G218gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT21), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n413_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n409_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n418_), .A2(KEYINPUT84), .B1(new_n406_), .B2(new_n405_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n408_), .A2(new_n420_), .A3(new_n409_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n415_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  OAI221_X1 g221(.A(new_n415_), .B1(new_n408_), .B2(new_n409_), .C1(new_n406_), .C2(new_n405_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n414_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n417_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G183gat), .A2(G190gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT23), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT23), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G183gat), .A3(G190gat), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n426_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(G169gat), .A2(G176gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT25), .B(G183gat), .Z(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT26), .B(G190gat), .Z(new_n435_));
  OAI221_X1 g234(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n429_), .B2(new_n427_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n429_), .B2(new_n427_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT74), .B(G176gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT22), .B(G169gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n432_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n404_), .B1(new_n425_), .B2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n436_), .A2(new_n443_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n446_), .B(new_n417_), .C1(new_n422_), .C2(new_n424_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G226gat), .A2(G233gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n450_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n403_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n403_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n392_), .A2(new_n391_), .A3(new_n386_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT93), .B1(new_n357_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n387_), .A2(new_n358_), .A3(new_n389_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n354_), .B(new_n355_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT93), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n458_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT33), .B(new_n357_), .C1(new_n390_), .C2(new_n393_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n454_), .A2(new_n457_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n390_), .A2(new_n357_), .A3(new_n393_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n394_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n452_), .A2(new_n453_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n456_), .A2(KEYINPUT32), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n470_), .A2(new_n471_), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n398_), .A2(new_n467_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G228gat), .ZN(new_n476_));
  INV_X1    g275(.A(G233gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT82), .B1(new_n380_), .B2(KEYINPUT29), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n425_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n479_), .A3(new_n425_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n485_), .A2(KEYINPUT81), .ZN(new_n486_));
  INV_X1    g285(.A(new_n483_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n484_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(new_n481_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G22gat), .B(G50gat), .Z(new_n490_));
  INV_X1    g289(.A(KEYINPUT28), .ZN(new_n491_));
  INV_X1    g290(.A(new_n380_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n380_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT80), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT28), .B1(new_n380_), .B2(KEYINPUT29), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n490_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT80), .B1(new_n494_), .B2(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n490_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n486_), .A2(new_n489_), .A3(new_n501_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n505_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n489_), .A2(new_n485_), .A3(KEYINPUT81), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n454_), .A2(new_n457_), .A3(KEYINPUT27), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT27), .B1(new_n454_), .B2(new_n457_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n469_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n475_), .A2(new_n511_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT75), .B(KEYINPUT76), .Z(new_n517_));
  NAND2_X1  g316(.A1(G227gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G15gat), .B(G43gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G71gat), .B(G99gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n519_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(KEYINPUT77), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(KEYINPUT77), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n526_), .B2(new_n523_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n383_), .B(KEYINPUT31), .Z(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT94), .B1(new_n516_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n469_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n514_), .A2(KEYINPUT95), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n514_), .A2(KEYINPUT95), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n535_), .B(new_n511_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539_));
  INV_X1    g338(.A(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n394_), .A2(new_n395_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n394_), .A2(KEYINPUT92), .A3(new_n395_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  AND4_X1   g344(.A1(new_n457_), .A2(new_n454_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n468_), .A2(new_n394_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n474_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n510_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n507_), .A2(new_n508_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n507_), .A2(new_n508_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n533_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n454_), .A2(new_n457_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT27), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n454_), .A2(new_n457_), .A3(KEYINPUT27), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n539_), .B(new_n540_), .C1(new_n551_), .C2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n532_), .A2(new_n538_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT67), .ZN(new_n564_));
  XOR2_X1   g363(.A(G134gat), .B(G162gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n335_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n320_), .A2(new_n242_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n572_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n573_), .A2(new_n579_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(KEYINPUT68), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n567_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n578_), .A2(new_n588_), .A3(new_n566_), .A4(new_n580_), .ZN(new_n589_));
  OAI211_X1 g388(.A(KEYINPUT69), .B(new_n567_), .C1(new_n582_), .C2(new_n584_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n562_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n350_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n533_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT97), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n562_), .A2(new_n268_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n581_), .A2(new_n567_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(KEYINPUT37), .A3(new_n589_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n591_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n237_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(new_n348_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n203_), .A3(new_n469_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n595_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT98), .ZN(G1324gat));
  NOR2_X1   g411(.A1(new_n536_), .A2(new_n537_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n593_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT39), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n606_), .A2(new_n204_), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g418(.A(G15gat), .B1(new_n593_), .B2(new_n540_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT41), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n605_), .A2(G15gat), .A3(new_n540_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1326gat));
  OAI21_X1  g422(.A(G22gat), .B1(new_n593_), .B2(new_n511_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT42), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n511_), .A2(G22gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n605_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT99), .Z(G1327gat));
  NAND3_X1  g427(.A1(new_n603_), .A2(new_n268_), .A3(new_n348_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n561_), .A2(new_n538_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n545_), .A2(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n631_));
  OAI22_X1  g430(.A1(new_n631_), .A2(new_n510_), .B1(new_n559_), .B2(new_n554_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n539_), .B1(new_n632_), .B2(new_n540_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n602_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT43), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n636_), .B(new_n602_), .C1(new_n630_), .C2(new_n633_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n629_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT100), .B1(new_n638_), .B2(KEYINPUT44), .ZN(new_n639_));
  INV_X1    g438(.A(new_n629_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n637_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n562_), .B2(new_n602_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n639_), .A2(new_n646_), .B1(KEYINPUT44), .B2(new_n638_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n469_), .ZN(new_n648_));
  INV_X1    g447(.A(G29gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n591_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n603_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n348_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n596_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n469_), .A2(new_n649_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT101), .ZN(new_n656_));
  OAI22_X1  g455(.A1(new_n648_), .A2(new_n649_), .B1(new_n654_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(new_n654_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n614_), .A2(G36gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT45), .B1(new_n654_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT44), .B(new_n640_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n613_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n639_), .B2(new_n646_), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT102), .B(KEYINPUT46), .Z(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(KEYINPUT103), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT103), .B1(new_n669_), .B2(new_n670_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n661_), .A2(new_n663_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n614_), .B1(new_n638_), .B2(KEYINPUT44), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n638_), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n644_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n678_), .B2(G36gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n673_), .B1(new_n679_), .B2(KEYINPUT46), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT46), .B(new_n664_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(KEYINPUT104), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n671_), .A2(new_n672_), .B1(new_n680_), .B2(new_n682_), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n647_), .A2(G43gat), .A3(new_n531_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G43gat), .B1(new_n658_), .B2(new_n531_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g487(.A(G50gat), .B1(new_n658_), .B2(new_n510_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n510_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n647_), .B2(new_n690_), .ZN(G1331gat));
  NAND2_X1  g490(.A1(new_n604_), .A2(new_n652_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT105), .Z(new_n693_));
  AND2_X1   g492(.A1(new_n562_), .A2(new_n267_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n219_), .A3(new_n469_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n592_), .A2(new_n237_), .A3(new_n267_), .A4(new_n652_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT106), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n469_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n219_), .ZN(G1332gat));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n217_), .A3(new_n613_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n613_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(G64gat), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1333gat));
  INV_X1    g505(.A(G71gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n698_), .B2(new_n531_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT49), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n695_), .A2(new_n707_), .A3(new_n531_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1334gat));
  INV_X1    g510(.A(G78gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n698_), .B2(new_n510_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT50), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n695_), .A2(new_n712_), .A3(new_n510_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1335gat));
  NAND4_X1  g515(.A1(new_n694_), .A2(new_n650_), .A3(new_n603_), .A4(new_n652_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n469_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n635_), .A2(new_n637_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n237_), .A2(new_n268_), .A3(new_n348_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT108), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT109), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n469_), .A2(G85gat), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT110), .Z(new_n726_));
  AOI21_X1  g525(.A(new_n719_), .B1(new_n724_), .B2(new_n726_), .ZN(G1336gat));
  NAND3_X1  g526(.A1(new_n718_), .A2(new_n279_), .A3(new_n613_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n724_), .A2(new_n613_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n279_), .ZN(G1337gat));
  NAND4_X1  g529(.A1(new_n718_), .A2(new_n531_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G99gat), .B1(new_n723_), .B2(new_n540_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n275_), .A3(new_n510_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G106gat), .B1(new_n723_), .B2(new_n511_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT52), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT52), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g539(.A1(new_n268_), .A2(new_n345_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n334_), .A2(new_n337_), .A3(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n321_), .A2(new_n322_), .A3(KEYINPUT55), .A4(new_n331_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT113), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n336_), .A2(new_n746_), .A3(KEYINPUT55), .A4(new_n322_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n310_), .A2(new_n336_), .A3(KEYINPUT111), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n321_), .A2(new_n302_), .A3(new_n309_), .A4(new_n331_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n315_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n743_), .B(new_n748_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT112), .B(new_n315_), .C1(new_n749_), .C2(new_n752_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n342_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT56), .B(new_n342_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n741_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n252_), .A2(new_n249_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n247_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n264_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n266_), .A2(new_n764_), .A3(KEYINPUT114), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n266_), .A2(new_n764_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n343_), .A2(new_n345_), .B1(new_n765_), .B2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT57), .B(new_n591_), .C1(new_n761_), .C2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n765_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n345_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n345_), .A3(KEYINPUT115), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n760_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT111), .B1(new_n310_), .B2(new_n336_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n750_), .A2(new_n751_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n316_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT112), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n743_), .A2(new_n748_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n753_), .A2(new_n754_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n342_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n776_), .B1(new_n777_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n601_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n776_), .B(KEYINPUT58), .C1(new_n777_), .C2(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n591_), .B1(new_n761_), .B2(new_n769_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n770_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n788_), .A2(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT119), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n603_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n601_), .A2(new_n237_), .A3(new_n348_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n268_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n613_), .A2(new_n510_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n469_), .A3(new_n531_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(G113gat), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n267_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n786_), .A2(new_n787_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n811_), .A2(KEYINPUT116), .A3(new_n602_), .A4(new_n789_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n793_), .A3(new_n770_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n788_), .B2(new_n789_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n603_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n815_), .A2(new_n803_), .A3(KEYINPUT117), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n815_), .B2(new_n803_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n806_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n808_), .B(new_n810_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n803_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n815_), .A2(new_n803_), .A3(KEYINPUT117), .ZN(new_n824_));
  INV_X1    g623(.A(new_n806_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n268_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n826_), .A2(KEYINPUT118), .A3(new_n809_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT118), .B1(new_n826_), .B2(new_n809_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n820_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT120), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n820_), .B(new_n831_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1340gat));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n348_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n818_), .B(new_n835_), .C1(KEYINPUT60), .C2(new_n834_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n808_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n818_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n348_), .B(new_n837_), .C1(new_n838_), .C2(KEYINPUT59), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n839_), .B2(new_n834_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n818_), .A2(new_n841_), .A3(new_n237_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n603_), .B(new_n837_), .C1(new_n838_), .C2(KEYINPUT59), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n841_), .ZN(G1342gat));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n838_), .B2(new_n591_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT121), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(new_n845_), .C1(new_n838_), .C2(new_n591_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n837_), .B1(new_n838_), .B2(KEYINPUT59), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n601_), .A2(new_n845_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT122), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n847_), .A2(new_n849_), .B1(new_n850_), .B2(new_n852_), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n823_), .A2(new_n824_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n540_), .A2(new_n469_), .A3(new_n510_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n854_), .A2(new_n613_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n268_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT123), .B(G141gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n652_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n237_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1346gat));
  INV_X1    g663(.A(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G162gat), .B1(new_n865_), .B2(new_n601_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n591_), .A2(G162gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n865_), .B2(new_n867_), .ZN(G1347gat));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n614_), .A2(new_n510_), .A3(new_n534_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n804_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n267_), .ZN(new_n872_));
  INV_X1    g671(.A(G169gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n441_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT62), .B(G169gat), .C1(new_n871_), .C2(new_n267_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(G1348gat));
  INV_X1    g676(.A(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n652_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n854_), .A2(new_n510_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n614_), .A2(new_n534_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n881_), .A2(G176gat), .A3(new_n652_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n879_), .A2(new_n440_), .B1(new_n880_), .B2(new_n882_), .ZN(G1349gat));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n237_), .A3(new_n881_), .ZN(new_n884_));
  INV_X1    g683(.A(G183gat), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n237_), .A2(new_n434_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n885_), .B1(new_n878_), .B2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n871_), .B2(new_n601_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n591_), .A2(new_n435_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n871_), .B2(new_n889_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n614_), .A2(new_n531_), .A3(new_n554_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n823_), .A2(new_n824_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT124), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n823_), .A2(new_n894_), .A3(new_n824_), .A4(new_n891_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n267_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n406_), .ZN(G1352gat));
  AOI21_X1  g696(.A(new_n348_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(G204gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n405_), .B2(new_n898_), .ZN(G1353gat));
  AOI21_X1  g699(.A(new_n603_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n816_), .A2(new_n817_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n894_), .B1(new_n902_), .B2(new_n891_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n895_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT125), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n907_), .B(KEYINPUT126), .Z(new_n908_));
  OAI211_X1 g707(.A(new_n905_), .B(new_n908_), .C1(KEYINPUT125), .C2(new_n906_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n908_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n901_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n906_), .A2(KEYINPUT125), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n909_), .A2(new_n914_), .ZN(G1354gat));
  NAND2_X1  g714(.A1(new_n602_), .A2(G218gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n591_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n650_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n917_), .B1(new_n920_), .B2(new_n922_), .ZN(G1355gat));
endmodule


