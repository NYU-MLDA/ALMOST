//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G1gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT71), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT71), .A2(G8gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n203_), .A2(new_n205_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT72), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n204_), .A2(G1gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n202_), .A2(KEYINPUT70), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT71), .A2(G8gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(KEYINPUT71), .A2(G8gat), .ZN(new_n216_));
  OAI22_X1  g015(.A1(new_n213_), .A2(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT72), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT14), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(G15gat), .B(G22gat), .Z(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT73), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n224_));
  AOI211_X1 g023(.A(new_n224_), .B(new_n221_), .C1(new_n212_), .C2(new_n219_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G1gat), .B(G8gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n223_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n210_), .A2(KEYINPUT72), .A3(new_n211_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n218_), .B1(new_n217_), .B2(KEYINPUT14), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n222_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n224_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n220_), .A2(KEYINPUT73), .A3(new_n222_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n226_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(G231gat), .B(G233gat), .C1(new_n228_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(G71gat), .ZN(new_n237_));
  INV_X1    g036(.A(G71gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(KEYINPUT65), .ZN(new_n239_));
  OAI21_X1  g038(.A(G78gat), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(KEYINPUT65), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(G71gat), .ZN(new_n242_));
  INV_X1    g041(.A(G78gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G57gat), .ZN(new_n246_));
  INV_X1    g045(.A(G57gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G64gat), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT11), .B1(new_n246_), .B2(new_n248_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n240_), .B(new_n244_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n243_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n227_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n232_), .A2(new_n233_), .A3(new_n226_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G231gat), .A2(G233gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n235_), .A2(new_n256_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G127gat), .B(G155gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G183gat), .B(G211gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT17), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(KEYINPUT74), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n256_), .B1(new_n235_), .B2(new_n260_), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n262_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n267_), .A2(KEYINPUT17), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n270_), .B(new_n273_), .C1(new_n262_), .C2(new_n271_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT37), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT37), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G29gat), .B(G36gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G43gat), .B(G50gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n279_), .B(KEYINPUT68), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT15), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n286_), .A3(KEYINPUT15), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT64), .B(G92gat), .Z(new_n292_));
  INV_X1    g091(.A(KEYINPUT9), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(G85gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G85gat), .B(G92gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT9), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT10), .B(G99gat), .Z(new_n298_));
  INV_X1    g097(.A(G106gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G99gat), .A2(G106gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT6), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G99gat), .A3(G106gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n294_), .A2(new_n297_), .A3(new_n300_), .A4(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT7), .ZN(new_n307_));
  INV_X1    g106(.A(G99gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(new_n299_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI211_X1 g110(.A(KEYINPUT8), .B(new_n295_), .C1(new_n311_), .C2(new_n305_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT8), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n305_), .A2(new_n310_), .A3(new_n309_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n296_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n306_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n291_), .A2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n316_), .A2(new_n287_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G232gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT34), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT35), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n318_), .A3(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n321_), .A2(new_n322_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G190gat), .B(G218gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G134gat), .B(G162gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT36), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n325_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n327_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n330_), .B(KEYINPUT36), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n277_), .B(new_n278_), .C1(new_n333_), .C2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n332_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n334_), .B1(new_n338_), .B2(new_n326_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n327_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n276_), .A4(KEYINPUT37), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n275_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G230gat), .A2(G233gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n316_), .A2(new_n256_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n302_), .A2(new_n304_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n309_), .A2(new_n310_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n296_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT8), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n314_), .A2(new_n313_), .A3(new_n296_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n251_), .A2(new_n255_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n306_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n345_), .B1(new_n346_), .B2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT66), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(KEYINPUT67), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n316_), .A2(new_n256_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n352_), .B2(new_n306_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(KEYINPUT67), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n346_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n345_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n355_), .A2(KEYINPUT66), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n356_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G120gat), .B(G148gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT5), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G176gat), .B(G204gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n370_), .B(new_n371_), .Z(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n372_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n356_), .A2(new_n366_), .A3(new_n367_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT13), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(KEYINPUT13), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n344_), .A2(KEYINPUT77), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  INV_X1    g181(.A(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT23), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT25), .B(G183gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT26), .B(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT24), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(G169gat), .B2(G176gat), .ZN(new_n398_));
  INV_X1    g197(.A(G169gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n386_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n395_), .A2(new_n396_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n386_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n392_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n394_), .A2(KEYINPUT79), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT79), .B1(new_n394_), .B2(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n384_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT80), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G113gat), .B(G120gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n394_), .A2(new_n403_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n384_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n404_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n407_), .A2(new_n412_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(G15gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT30), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n412_), .B1(new_n407_), .B2(new_n417_), .ZN(new_n425_));
  OR3_X1    g224(.A1(new_n419_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G155gat), .A2(G162gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n433_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(G155gat), .ZN(new_n435_));
  INV_X1    g234(.A(G162gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT1), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n431_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n429_), .B(KEYINPUT3), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT2), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n437_), .A3(new_n432_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT29), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G228gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G211gat), .B(G218gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT85), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT21), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G197gat), .B(G204gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G197gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n456_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT21), .B(new_n459_), .C1(new_n460_), .C2(KEYINPUT84), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n457_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n456_), .A2(new_n455_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n454_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n448_), .A2(KEYINPUT83), .A3(KEYINPUT29), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n451_), .A2(new_n452_), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n449_), .A2(new_n465_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469_));
  INV_X1    g268(.A(new_n452_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n457_), .A2(new_n461_), .B1(new_n454_), .B2(new_n463_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(KEYINPUT29), .B2(new_n448_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT86), .B1(new_n473_), .B2(new_n452_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n467_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT28), .B1(new_n448_), .B2(KEYINPUT29), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n440_), .B(KEYINPUT82), .ZN(new_n477_));
  INV_X1    g276(.A(new_n447_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT28), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT29), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G22gat), .B(G50gat), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n476_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G78gat), .B(G106gat), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n467_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n484_), .A2(new_n485_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n487_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT87), .B1(new_n490_), .B2(new_n491_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n428_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n492_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n493_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n428_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n494_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n472_), .B1(new_n415_), .B2(new_n404_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT88), .B1(new_n387_), .B2(new_n390_), .ZN(new_n505_));
  OR2_X1    g304(.A1(G183gat), .A2(G190gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n392_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n387_), .A2(KEYINPUT88), .A3(new_n390_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n403_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n465_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT19), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n504_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n513_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n415_), .A2(new_n472_), .A3(new_n404_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n465_), .B2(new_n510_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n515_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G8gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT18), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G64gat), .B(G92gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n514_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT95), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n516_), .A2(new_n518_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n513_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n510_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n517_), .B1(new_n529_), .B2(new_n472_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n465_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n515_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n523_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n523_), .B(KEYINPUT94), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n515_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n516_), .A2(new_n518_), .A3(new_n515_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n526_), .A2(KEYINPUT27), .A3(new_n535_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT27), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n523_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n525_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n479_), .A2(new_n412_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n448_), .A2(new_n411_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(KEYINPUT4), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G225gat), .A2(G233gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT4), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n448_), .A2(new_n550_), .A3(new_n411_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n448_), .B(new_n412_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n548_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G1gat), .B(G29gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G85gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT0), .B(G57gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n552_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n544_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n565_));
  INV_X1    g364(.A(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n523_), .A2(KEYINPUT32), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n528_), .A2(new_n532_), .A3(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n565_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n563_), .A2(KEYINPUT93), .A3(new_n570_), .A4(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n553_), .A2(new_n549_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n560_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT91), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n547_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n581_), .A3(new_n560_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n576_), .A2(new_n579_), .A3(new_n580_), .A4(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(KEYINPUT90), .A2(KEYINPUT33), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n562_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n525_), .A2(new_n542_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n583_), .B(new_n585_), .C1(new_n586_), .C2(KEYINPUT89), .ZN(new_n587_));
  INV_X1    g386(.A(new_n542_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n533_), .A3(KEYINPUT89), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n562_), .A2(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n572_), .B(new_n573_), .C1(new_n587_), .C2(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n495_), .A2(new_n501_), .A3(new_n496_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n503_), .A2(new_n564_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n257_), .A2(new_n258_), .A3(new_n287_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n287_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n287_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n257_), .A2(new_n291_), .A3(new_n258_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n595_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G113gat), .B(G141gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G169gat), .B(G197gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  AND3_X1   g405(.A1(new_n599_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n594_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT77), .B1(new_n344_), .B2(new_n380_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n381_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT96), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n381_), .A2(new_n610_), .A3(new_n611_), .A4(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n563_), .B(KEYINPUT97), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n617_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(KEYINPUT98), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n615_), .A3(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n619_), .A2(KEYINPUT38), .A3(new_n622_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n333_), .A2(new_n336_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n594_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n275_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n380_), .A2(new_n609_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n566_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT99), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n625_), .A2(new_n626_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n208_), .A2(new_n209_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n616_), .A2(new_n637_), .A3(new_n544_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n628_), .A2(new_n544_), .A3(new_n630_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(KEYINPUT100), .A2(KEYINPUT39), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n207_), .B1(KEYINPUT100), .B2(KEYINPUT39), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n641_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n635_), .B1(new_n639_), .B2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n638_), .B(KEYINPUT40), .C1(new_n645_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  OAI21_X1  g448(.A(G15gat), .B1(new_n631_), .B2(new_n428_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT41), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n612_), .A2(G15gat), .A3(new_n428_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n495_), .A2(new_n496_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G22gat), .B1(new_n631_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n654_), .A2(G22gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n612_), .B2(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(new_n380_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n594_), .A2(new_n609_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n563_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n337_), .A2(new_n341_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n594_), .B2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n495_), .A2(new_n496_), .A3(new_n428_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n501_), .B1(new_n500_), .B2(new_n494_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n564_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n592_), .A2(new_n593_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n664_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n666_), .A2(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n380_), .A2(new_n609_), .A3(new_n275_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(KEYINPUT44), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n674_), .B2(new_n675_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n617_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(G29gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n663_), .B1(new_n678_), .B2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(G36gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n662_), .A2(new_n682_), .A3(new_n544_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  INV_X1    g483(.A(new_n544_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n676_), .A2(new_n677_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(new_n682_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(KEYINPUT46), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n687_), .B(new_n689_), .ZN(G1329gat));
  AOI21_X1  g489(.A(G43gat), .B1(new_n662_), .B2(new_n501_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n428_), .A2(new_n383_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n678_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g493(.A1(new_n654_), .A2(G50gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT103), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n662_), .A2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n676_), .A2(new_n677_), .A3(new_n654_), .ZN(new_n698_));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n698_), .B2(new_n699_), .ZN(G1331gat));
  NAND4_X1  g499(.A1(new_n628_), .A2(new_n609_), .A3(new_n275_), .A4(new_n380_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n701_), .A2(new_n247_), .A3(new_n566_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n609_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n594_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n344_), .A2(new_n660_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n707_), .A2(KEYINPUT104), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(KEYINPUT104), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n679_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n702_), .B1(new_n710_), .B2(new_n247_), .ZN(G1332gat));
  OAI21_X1  g510(.A(G64gat), .B1(new_n701_), .B2(new_n685_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT48), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n245_), .A3(new_n544_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n701_), .B2(new_n428_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n707_), .A2(new_n238_), .A3(new_n501_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n701_), .B2(new_n654_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  INV_X1    g520(.A(new_n654_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n707_), .A2(new_n243_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1335gat));
  NAND3_X1  g523(.A1(new_n380_), .A2(new_n609_), .A3(new_n629_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n666_), .B2(new_n673_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(G85gat), .A3(new_n563_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n704_), .A2(new_n627_), .A3(new_n629_), .A4(new_n380_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT105), .ZN(new_n729_));
  AOI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n679_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT106), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT106), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g532(.A(G92gat), .B1(new_n729_), .B2(new_n544_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n544_), .A2(new_n292_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n726_), .B2(new_n735_), .ZN(G1337gat));
  AOI21_X1  g535(.A(new_n308_), .B1(new_n726_), .B2(new_n501_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n501_), .A2(new_n298_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n729_), .A2(new_n740_), .B1(KEYINPUT108), .B2(KEYINPUT51), .ZN(new_n741_));
  OR2_X1    g540(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n739_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n729_), .A2(new_n299_), .A3(new_n722_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n725_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n672_), .B1(new_n671_), .B2(new_n664_), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT43), .B(new_n665_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n722_), .B(new_n747_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT109), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n654_), .B(new_n725_), .C1(new_n666_), .C2(new_n673_), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT110), .B(KEYINPUT52), .C1(new_n754_), .C2(new_n299_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n750_), .A2(new_n757_), .A3(new_n751_), .A4(G106gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(KEYINPUT110), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n746_), .B1(new_n756_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n746_), .B(new_n762_), .C1(new_n756_), .C2(new_n760_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1339gat));
  AOI21_X1  g565(.A(new_n358_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n362_), .B1(new_n346_), .B2(new_n354_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n345_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(KEYINPUT55), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n361_), .A2(KEYINPUT55), .A3(new_n365_), .A4(new_n345_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n372_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT117), .A3(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT56), .B(new_n372_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n345_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n366_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n374_), .B1(new_n784_), .B2(new_n773_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n785_), .B2(KEYINPUT56), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n777_), .A2(new_n780_), .A3(new_n786_), .A4(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n606_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(KEYINPUT115), .A3(new_n790_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n601_), .A2(new_n596_), .A3(new_n602_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n607_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n375_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n664_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT58), .B1(new_n788_), .B2(new_n798_), .ZN(new_n801_));
  AOI211_X1 g600(.A(KEYINPUT113), .B(new_n374_), .C1(new_n784_), .C2(new_n773_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n776_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n375_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT112), .B(new_n375_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n803_), .A2(new_n776_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n775_), .B1(KEYINPUT113), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n804_), .A2(new_n807_), .A3(new_n808_), .A4(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n796_), .A2(new_n797_), .A3(new_n376_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n627_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n800_), .A2(new_n801_), .B1(new_n813_), .B2(KEYINPUT57), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n813_), .A2(KEYINPUT57), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n629_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n378_), .A2(new_n609_), .A3(new_n379_), .ZN(new_n817_));
  OR3_X1    g616(.A1(new_n817_), .A2(new_n342_), .A3(KEYINPUT54), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n817_), .B2(new_n342_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n617_), .A2(new_n544_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n667_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT118), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n825_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n609_), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n828_), .A2(G113gat), .A3(new_n609_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1340gat));
  OAI21_X1  g633(.A(G120gat), .B1(new_n831_), .B2(new_n660_), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n660_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(KEYINPUT60), .B2(new_n836_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n828_), .B2(new_n838_), .ZN(G1341gat));
  AOI21_X1  g638(.A(G127gat), .B1(new_n826_), .B2(new_n275_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n275_), .A2(G127gat), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT119), .Z(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT120), .B(new_n841_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n847_), .ZN(G1342gat));
  XNOR2_X1  g647(.A(KEYINPUT121), .B(G134gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n831_), .A2(new_n665_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G134gat), .B1(new_n826_), .B2(new_n627_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n811_), .A2(new_n812_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n627_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n813_), .A2(KEYINPUT57), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n788_), .A2(new_n798_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n664_), .A3(new_n799_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n858_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n820_), .B1(new_n863_), .B2(new_n629_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n497_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n823_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n703_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n380_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n866_), .A2(new_n629_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n866_), .B2(new_n665_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n627_), .A2(new_n436_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n866_), .B2(new_n876_), .ZN(G1347gat));
  NOR3_X1   g676(.A1(new_n679_), .A2(new_n685_), .A3(new_n502_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n703_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n864_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  INV_X1    g680(.A(new_n879_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n822_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n883_), .A3(G169gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT62), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n399_), .A2(KEYINPUT62), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n880_), .A2(new_n883_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n880_), .A2(new_n883_), .A3(new_n892_), .A4(new_n889_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n887_), .A2(new_n888_), .A3(new_n891_), .A4(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n822_), .A2(new_n385_), .A3(new_n882_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1348gat));
  NAND2_X1  g695(.A1(new_n822_), .A2(new_n878_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n660_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n386_), .ZN(G1349gat));
  OR3_X1    g698(.A1(new_n897_), .A2(new_n395_), .A3(new_n629_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n629_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(G183gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n903_), .B2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n897_), .B2(new_n665_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n627_), .A2(new_n396_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n897_), .B2(new_n907_), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n685_), .A2(new_n563_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n865_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n910_), .B(new_n703_), .C1(KEYINPUT126), .C2(G197gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT126), .B(G197gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n865_), .A2(new_n909_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n609_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n911_), .A2(new_n914_), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n380_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g716(.A(KEYINPUT63), .B(G211gat), .Z(new_n918_));
  NAND3_X1  g717(.A1(new_n910_), .A2(new_n275_), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(KEYINPUT127), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n913_), .B2(new_n629_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n919_), .A2(KEYINPUT127), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1354gat));
  OR3_X1    g724(.A1(new_n913_), .A2(G218gat), .A3(new_n854_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G218gat), .B1(new_n913_), .B2(new_n665_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1355gat));
endmodule


