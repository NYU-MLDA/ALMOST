//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(KEYINPUT93), .A2(KEYINPUT2), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT93), .A2(KEYINPUT2), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT94), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT94), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n208_), .B(new_n203_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n209_));
  OR4_X1    g008(.A1(KEYINPUT92), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n210_));
  OAI22_X1  g009(.A1(KEYINPUT92), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n207_), .A2(new_n209_), .A3(new_n210_), .A4(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT91), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n217_), .B(KEYINPUT1), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n216_), .ZN(new_n220_));
  INV_X1    g019(.A(G141gat), .ZN(new_n221_));
  INV_X1    g020(.A(G148gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n203_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n202_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G218gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(G211gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT97), .ZN(new_n228_));
  INV_X1    g027(.A(G211gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(G218gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  AOI211_X1 g031(.A(new_n227_), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(new_n232_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n225_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT96), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(KEYINPUT96), .A2(G233gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(G228gat), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT98), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT98), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n242_), .B(new_n243_), .C1(new_n225_), .C2(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n235_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n218_), .A2(new_n224_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT95), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT95), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n218_), .A2(new_n249_), .A3(new_n224_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n246_), .B(new_n240_), .C1(new_n251_), .C2(new_n202_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT100), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT100), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n245_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G22gat), .B(G50gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n258_));
  INV_X1    g057(.A(new_n250_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n249_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n258_), .B(new_n202_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n251_), .B2(new_n202_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n259_), .A2(new_n260_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT28), .B1(new_n265_), .B2(KEYINPUT29), .ZN(new_n266_));
  INV_X1    g065(.A(new_n257_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n261_), .A3(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G78gat), .B(G106gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n264_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(KEYINPUT99), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n264_), .B2(new_n268_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n254_), .B(new_n256_), .C1(new_n271_), .C2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n254_), .A2(new_n256_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G226gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT19), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT86), .B(G176gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT84), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G183gat), .ZN(new_n288_));
  INV_X1    g087(.A(G190gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT23), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  OR3_X1    g091(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT23), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(new_n289_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n287_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G183gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n288_), .A2(KEYINPUT25), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n289_), .A2(KEYINPUT26), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n297_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n293_), .A2(new_n290_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n285_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n306_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n296_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n235_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n297_), .B1(new_n286_), .B2(new_n309_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n299_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT83), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n302_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(KEYINPUT81), .B(G183gat), .Z(new_n321_));
  OAI221_X1 g120(.A(new_n304_), .B1(new_n315_), .B2(new_n299_), .C1(new_n321_), .C2(new_n298_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n294_), .B(new_n314_), .C1(new_n320_), .C2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n307_), .B1(new_n321_), .B2(G190gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT87), .B1(new_n282_), .B2(new_n283_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n282_), .A2(KEYINPUT87), .A3(new_n283_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n324_), .B(new_n286_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(new_n246_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n281_), .B1(new_n313_), .B2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G8gat), .B(G36gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT20), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n312_), .B2(new_n235_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n281_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n328_), .A2(new_n246_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n330_), .A2(new_n336_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n340_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n281_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n296_), .A2(new_n311_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n337_), .B1(new_n345_), .B2(new_n246_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n329_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n339_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n336_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT103), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n342_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n313_), .A2(new_n329_), .A3(new_n281_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n339_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n354_), .A2(KEYINPUT103), .A3(new_n336_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT27), .B1(new_n351_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n330_), .A2(new_n341_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n335_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n342_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT27), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n279_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT89), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n363_), .B(new_n365_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(KEYINPUT89), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT90), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT102), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n247_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n368_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n370_), .A2(KEYINPUT102), .A3(new_n248_), .A4(new_n250_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n373_), .A2(KEYINPUT4), .A3(new_n375_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n371_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n373_), .A2(new_n378_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  AND3_X1   g186(.A1(new_n382_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n370_), .A2(KEYINPUT31), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n370_), .A2(KEYINPUT31), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT88), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n328_), .B(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G43gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n403_), .A3(new_n400_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n390_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n362_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n382_), .A2(KEYINPUT33), .A3(new_n383_), .A4(new_n387_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n378_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n377_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n387_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n373_), .A2(new_n411_), .A3(new_n375_), .A4(new_n376_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n359_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n376_), .A2(new_n375_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT102), .B1(new_n265_), .B2(new_n370_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n377_), .A2(new_n381_), .B1(new_n421_), .B2(new_n378_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT33), .B1(new_n422_), .B2(new_n387_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n418_), .A2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n336_), .A2(KEYINPUT32), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n354_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n330_), .B2(new_n341_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n389_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n382_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n279_), .B1(new_n424_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n274_), .A2(new_n278_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n361_), .A2(new_n433_), .A3(new_n390_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n407_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n409_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G169gat), .B(G197gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  XNOR2_X1  g239(.A(G29gat), .B(G36gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT69), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT69), .ZN(new_n443_));
  INV_X1    g242(.A(G29gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(G36gat), .ZN(new_n445_));
  INV_X1    g244(.A(G36gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(G29gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n443_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G43gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(G50gat), .ZN(new_n451_));
  INV_X1    g250(.A(G50gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(G43gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT70), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(G43gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(G50gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n449_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n442_), .A2(new_n448_), .A3(new_n454_), .A4(new_n458_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n466_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n460_), .A2(new_n467_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G229gat), .A2(G233gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n465_), .B(new_n466_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT15), .ZN(new_n476_));
  AND4_X1   g275(.A1(new_n442_), .A2(new_n448_), .A3(new_n454_), .A4(new_n458_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n442_), .A2(new_n448_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n460_), .A2(new_n468_), .A3(KEYINPUT15), .ZN(new_n480_));
  AOI211_X1 g279(.A(KEYINPUT77), .B(new_n475_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT77), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n474_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n473_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT76), .B1(new_n486_), .B2(new_n470_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n471_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(KEYINPUT76), .A3(new_n470_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n440_), .B1(new_n485_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n460_), .A2(new_n468_), .A3(KEYINPUT15), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT15), .B1(new_n460_), .B2(new_n468_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n474_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT77), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n483_), .A2(new_n482_), .A3(new_n474_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n486_), .A2(KEYINPUT76), .A3(new_n470_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(new_n487_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n499_), .A2(new_n473_), .B1(new_n501_), .B2(new_n489_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT78), .B1(new_n502_), .B2(new_n440_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n485_), .A2(new_n491_), .A3(KEYINPUT78), .A4(new_n440_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n493_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n485_), .A2(new_n491_), .A3(new_n440_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n504_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(KEYINPUT79), .A3(new_n493_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT80), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n437_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G85gat), .ZN(new_n517_));
  INV_X1    g316(.A(G92gat), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT9), .ZN(new_n519_));
  AND2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(KEYINPUT9), .B2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n524_));
  INV_X1    g323(.A(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT64), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT6), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n524_), .A2(new_n534_), .A3(new_n525_), .A4(new_n526_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n523_), .A2(new_n528_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G85gat), .B(G92gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  AOI211_X1 g342(.A(new_n537_), .B(new_n539_), .C1(new_n543_), .C2(new_n533_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n545_));
  INV_X1    g344(.A(G99gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n525_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n531_), .B1(G99gat), .B2(G106gat), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n529_), .A2(KEYINPUT6), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n540_), .B(new_n547_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n538_), .B1(new_n550_), .B2(new_n522_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n536_), .B1(new_n544_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n483_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT71), .Z(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT66), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n552_), .A2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT66), .B(new_n536_), .C1(new_n544_), .C2(new_n551_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n460_), .A2(new_n468_), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n563_), .A2(new_n564_), .B1(KEYINPUT35), .B2(new_n556_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n554_), .A2(new_n559_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n559_), .B1(new_n554_), .B2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G190gat), .B(G218gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT72), .ZN(new_n570_));
  XOR2_X1   g369(.A(G134gat), .B(G162gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT36), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n566_), .A2(new_n576_), .A3(new_n572_), .A4(new_n567_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n577_), .A2(new_n575_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT37), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n568_), .A2(KEYINPUT74), .A3(new_n573_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n577_), .A4(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT11), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT11), .ZN(new_n590_));
  INV_X1    g389(.A(G57gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(G64gat), .ZN(new_n592_));
  INV_X1    g391(.A(G64gat), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(G57gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n590_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n589_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n596_), .A3(KEYINPUT11), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n561_), .A2(new_n562_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n587_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n552_), .B(KEYINPUT12), .C1(new_n601_), .C2(new_n602_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n604_), .B(new_n608_), .C1(new_n606_), .C2(KEYINPUT12), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n587_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XOR2_X1   g411(.A(G176gat), .B(G204gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n610_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT13), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n603_), .B(new_n474_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT17), .B1(new_n619_), .B2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n619_), .B2(KEYINPUT75), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT17), .B(new_n623_), .C1(new_n619_), .C2(KEYINPUT75), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n586_), .A2(new_n616_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n516_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n390_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n462_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n361_), .A2(new_n433_), .A3(new_n390_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n430_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n387_), .B1(new_n421_), .B2(new_n411_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n359_), .B1(new_n640_), .B2(new_n413_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(new_n641_), .A3(new_n410_), .ZN(new_n642_));
  OAI22_X1  g441(.A1(new_n388_), .A2(new_n389_), .B1(new_n427_), .B2(new_n426_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n433_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n436_), .B1(new_n637_), .B2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n362_), .A2(new_n408_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n582_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n628_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n616_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n514_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n390_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n634_), .A2(new_n635_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n636_), .A2(new_n658_), .A3(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(new_n361_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n632_), .A2(new_n463_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n657_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n661_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n463_), .B1(new_n665_), .B2(KEYINPUT39), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n662_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n670_), .B(new_n671_), .Z(G1325gat));
  NAND2_X1  g471(.A1(new_n663_), .A2(new_n407_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(G15gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n673_), .B2(G15gat), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n632_), .A2(new_n395_), .A3(new_n407_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n657_), .B2(new_n279_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n279_), .A2(G22gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n631_), .B2(new_n685_), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n649_), .A2(new_n650_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n437_), .A2(new_n515_), .A3(new_n654_), .A4(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n444_), .A3(new_n633_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n586_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT107), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n693_), .B(KEYINPUT43), .C1(new_n437_), .C2(new_n586_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n580_), .A2(new_n585_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n407_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n691_), .B(new_n696_), .C1(new_n697_), .C2(new_n409_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT108), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n690_), .A2(new_n700_), .A3(new_n691_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n695_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n656_), .A2(new_n650_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n695_), .B2(new_n702_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n709_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n390_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(KEYINPUT110), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G29gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT110), .B1(new_n711_), .B2(new_n714_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n689_), .B1(new_n716_), .B2(new_n717_), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n688_), .A2(new_n446_), .A3(new_n661_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n661_), .B1(new_n709_), .B2(KEYINPUT44), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n446_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT46), .B(new_n720_), .C1(new_n722_), .C2(new_n446_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  NAND2_X1  g526(.A1(new_n712_), .A2(new_n713_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n436_), .A2(new_n450_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n710_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT109), .B1(new_n709_), .B2(KEYINPUT44), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n728_), .B(new_n729_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G43gat), .B1(new_n688_), .B2(new_n407_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT111), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n688_), .B2(new_n433_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n711_), .A2(new_n728_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n279_), .A2(new_n452_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  NAND3_X1  g542(.A1(new_n653_), .A2(new_n515_), .A3(new_n654_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n390_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n437_), .A2(new_n514_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n696_), .A2(new_n616_), .A3(new_n650_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n591_), .A3(new_n633_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n745_), .A2(new_n750_), .ZN(G1332gat));
  OAI21_X1  g550(.A(G64gat), .B1(new_n744_), .B2(new_n361_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT48), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n593_), .A3(new_n661_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n744_), .B2(new_n436_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT49), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n436_), .A2(G71gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n748_), .B2(new_n759_), .ZN(G1334gat));
  OAI21_X1  g559(.A(G78gat), .B1(new_n744_), .B2(new_n279_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT50), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n279_), .A2(G78gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n748_), .B2(new_n763_), .ZN(G1335gat));
  NAND3_X1  g563(.A1(new_n654_), .A2(new_n655_), .A3(new_n650_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n695_), .B2(new_n702_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n390_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n687_), .A2(new_n616_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n746_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n517_), .A3(new_n633_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n768_), .A2(new_n772_), .ZN(G1336gat));
  OAI21_X1  g572(.A(G92gat), .B1(new_n767_), .B2(new_n361_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n518_), .A3(new_n661_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1337gat));
  NAND2_X1  g575(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n407_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n770_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n766_), .A2(new_n407_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G99gat), .ZN(new_n781_));
  NOR2_X1   g580(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1338gat));
  AOI21_X1  g582(.A(new_n525_), .B1(new_n766_), .B2(new_n433_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT52), .B1(new_n784_), .B2(KEYINPUT114), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n279_), .B(new_n765_), .C1(new_n695_), .C2(new_n702_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n525_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n771_), .A2(new_n525_), .A3(new_n433_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(new_n525_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(KEYINPUT52), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n784_), .A2(KEYINPUT114), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n791_), .A3(KEYINPUT52), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n784_), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .A4(new_n790_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n793_), .A2(new_n798_), .ZN(G1339gat));
  XOR2_X1   g598(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n800_));
  NAND3_X1  g599(.A1(new_n630_), .A2(new_n515_), .A3(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n802_));
  INV_X1    g601(.A(new_n515_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n629_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT117), .B1(new_n609_), .B2(new_n587_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT55), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT117), .B(new_n809_), .C1(new_n609_), .C2(new_n587_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n609_), .A2(new_n587_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n614_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n614_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n610_), .A2(new_n614_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT79), .B1(new_n512_), .B2(new_n493_), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n507_), .B(new_n492_), .C1(new_n511_), .C2(new_n504_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT116), .B(new_n818_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n514_), .B2(new_n818_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n806_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(KEYINPUT118), .A3(new_n817_), .A4(new_n821_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n499_), .A2(new_n489_), .A3(new_n470_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n440_), .B1(new_n501_), .B2(new_n471_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n511_), .A2(new_n504_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n615_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n824_), .A2(new_n828_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n648_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT57), .A3(new_n648_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n818_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n815_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(KEYINPUT119), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(KEYINPUT119), .B2(new_n817_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n586_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n836_), .A2(new_n837_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n805_), .B1(new_n846_), .B2(new_n650_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n633_), .A2(new_n407_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n362_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n847_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n514_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n834_), .A2(new_n835_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n628_), .B1(new_n856_), .B2(new_n837_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT59), .B(new_n849_), .C1(new_n857_), .C2(new_n805_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n515_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n853_), .B1(new_n859_), .B2(new_n852_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n862_), .B(new_n853_), .C1(new_n859_), .C2(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1340gat));
  XOR2_X1   g663(.A(KEYINPUT122), .B(G120gat), .Z(new_n865_));
  OR2_X1    g664(.A1(new_n865_), .A2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n616_), .B2(KEYINPUT60), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n851_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n616_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n865_), .B2(new_n871_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n851_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n650_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n873_), .C1(new_n874_), .C2(new_n650_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n855_), .A2(new_n858_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n650_), .A2(new_n873_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n876_), .A2(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(G1342gat));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n851_), .A2(new_n882_), .A3(new_n649_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n586_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n882_), .ZN(G1343gat));
  INV_X1    g684(.A(new_n847_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n661_), .A2(new_n279_), .A3(new_n390_), .A4(new_n407_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n655_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT125), .B(G141gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1344gat));
  NOR2_X1   g690(.A1(new_n888_), .A2(new_n616_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n222_), .ZN(G1345gat));
  NOR2_X1   g692(.A1(new_n888_), .A2(new_n650_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT61), .B(G155gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n888_), .B2(new_n586_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n648_), .A2(G162gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n888_), .B2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n408_), .A2(new_n433_), .A3(new_n361_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n886_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n655_), .ZN(new_n903_));
  INV_X1    g702(.A(G169gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n900_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n283_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(G169gat), .C1(new_n902_), .C2(new_n655_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  NOR2_X1   g707(.A1(new_n902_), .A2(new_n616_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n282_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(G176gat), .B2(new_n909_), .ZN(G1349gat));
  NOR2_X1   g711(.A1(new_n902_), .A2(new_n650_), .ZN(new_n913_));
  MUX2_X1   g712(.A(new_n321_), .B(new_n301_), .S(new_n913_), .Z(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n902_), .B2(new_n586_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n649_), .A2(new_n305_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n902_), .B2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n436_), .A2(new_n433_), .A3(new_n390_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n361_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n886_), .A2(KEYINPUT127), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  INV_X1    g722(.A(new_n921_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n847_), .B2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n655_), .B1(new_n922_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(G197gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1352gat));
  AOI21_X1  g727(.A(new_n616_), .B1(new_n922_), .B2(new_n925_), .ZN(new_n929_));
  INV_X1    g728(.A(G204gat), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1353gat));
  XNOR2_X1  g730(.A(KEYINPUT63), .B(G211gat), .ZN(new_n932_));
  AOI211_X1 g731(.A(new_n650_), .B(new_n932_), .C1(new_n922_), .C2(new_n925_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n922_), .A2(new_n925_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n628_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  NAND3_X1  g736(.A1(new_n934_), .A2(new_n226_), .A3(new_n649_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n586_), .B1(new_n922_), .B2(new_n925_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n226_), .ZN(G1355gat));
endmodule


