//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n207_), .A3(new_n209_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n208_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT65), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n209_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT64), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n217_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n224_), .B2(new_n203_), .ZN(new_n225_));
  AOI211_X1 g024(.A(KEYINPUT8), .B(new_n202_), .C1(new_n223_), .C2(new_n209_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n213_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n230_), .B(new_n213_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G232gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT34), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(KEYINPUT35), .A3(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(KEYINPUT35), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n232_), .A2(new_n233_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(KEYINPUT69), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n239_), .A2(KEYINPUT69), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G190gat), .B(G218gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT67), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G134gat), .B(G162gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT36), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT68), .Z(new_n249_));
  AND2_X1   g048(.A1(new_n242_), .A2(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT70), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT70), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n246_), .B(KEYINPUT36), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(new_n241_), .A3(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(KEYINPUT37), .A3(new_n252_), .A4(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT37), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n240_), .A2(KEYINPUT71), .A3(new_n241_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT71), .B1(new_n240_), .B2(new_n241_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n253_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n260_), .B2(new_n250_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G1gat), .B(G8gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT72), .ZN(new_n264_));
  XOR2_X1   g063(.A(G15gat), .B(G22gat), .Z(new_n265_));
  NAND2_X1  g064(.A1(G1gat), .A2(G8gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(KEYINPUT14), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n264_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT73), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n268_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G57gat), .B(G64gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G71gat), .B(G78gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n275_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n271_), .B(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G127gat), .B(G155gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(G183gat), .B(G211gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT17), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n281_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n281_), .A2(new_n288_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n262_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT75), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G230gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n280_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n227_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n227_), .A2(new_n298_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT12), .A3(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(KEYINPUT12), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n297_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G120gat), .B(G148gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT5), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G176gat), .B(G204gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT66), .B(KEYINPUT13), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n313_), .B2(KEYINPUT13), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n295_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G204gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT89), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G204gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(G197gat), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT88), .B1(new_n323_), .B2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n318_), .A3(G197gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT21), .B1(new_n322_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n323_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G197gat), .A2(G204gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n330_), .A2(new_n331_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n333_), .A2(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT23), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n343_));
  INV_X1    g142(.A(G183gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(KEYINPUT23), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n342_), .A2(new_n343_), .B1(G190gat), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT26), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT78), .A3(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(KEYINPUT25), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT25), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G183gat), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .A4(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT79), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G169gat), .ZN(new_n358_));
  INV_X1    g157(.A(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT24), .A4(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n354_), .A2(new_n357_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G183gat), .A3(G190gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n340_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n369_), .B1(new_n373_), .B2(KEYINPUT81), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n375_), .B(new_n370_), .C1(new_n340_), .C2(new_n372_), .ZN(new_n376_));
  OAI22_X1  g175(.A1(new_n346_), .A2(new_n365_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n338_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n340_), .A2(new_n372_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n364_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT95), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n382_), .A3(new_n364_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT25), .B(G183gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n355_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n384_), .A2(new_n385_), .B1(new_n386_), .B2(new_n362_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n369_), .B1(new_n346_), .B2(new_n370_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(new_n334_), .A3(new_n389_), .A4(new_n337_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n378_), .A2(KEYINPUT20), .A3(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G8gat), .B(G36gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n388_), .A2(new_n389_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT96), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n402_), .A2(new_n338_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n402_), .B2(new_n338_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n338_), .B2(new_n377_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n394_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n395_), .B(new_n401_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT102), .B1(new_n407_), .B2(new_n408_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n405_), .A2(new_n406_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n402_), .A2(new_n338_), .A3(new_n403_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n391_), .A2(new_n394_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(KEYINPUT102), .B2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT27), .B(new_n409_), .C1(new_n416_), .C2(new_n401_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n408_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n391_), .A2(new_n394_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n400_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT98), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n409_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT27), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT98), .B(new_n400_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n417_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT82), .B(G15gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n377_), .B(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G71gat), .B(G99gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G43gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n431_), .B(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n435_), .A2(KEYINPUT83), .ZN(new_n436_));
  INV_X1    g235(.A(G134gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G127gat), .ZN(new_n438_));
  INV_X1    g237(.A(G127gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G134gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G120gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G113gat), .ZN(new_n443_));
  INV_X1    g242(.A(G113gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G120gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n438_), .A2(new_n440_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n449_), .B(KEYINPUT31), .Z(new_n450_));
  OR2_X1    g249(.A1(new_n436_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n435_), .A2(KEYINPUT83), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n436_), .A2(new_n452_), .A3(new_n450_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n455_));
  INV_X1    g254(.A(G141gat), .ZN(new_n456_));
  INV_X1    g255(.A(G148gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT85), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G155gat), .ZN(new_n469_));
  INV_X1    g268(.A(G162gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n465_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n464_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n456_), .A2(new_n457_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(KEYINPUT1), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n471_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n465_), .A2(KEYINPUT1), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n459_), .B(new_n475_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT29), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n338_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(G228gat), .A3(G233gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT90), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(KEYINPUT90), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n481_), .A2(KEYINPUT87), .B1(G228gat), .B2(G233gat), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(new_n338_), .C1(KEYINPUT87), .C2(new_n481_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G78gat), .B(G106gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT91), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT92), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .A4(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n480_), .A2(KEYINPUT29), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G22gat), .B(G50gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n493_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n491_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n501_), .A2(KEYINPUT93), .A3(new_n489_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT93), .B1(new_n501_), .B2(new_n489_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n490_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n491_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n506_), .A2(new_n507_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n449_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n480_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n474_), .A2(new_n449_), .A3(new_n479_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G225gat), .A2(G233gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n480_), .A2(new_n516_), .A3(new_n510_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n474_), .A2(new_n449_), .A3(new_n479_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n449_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n517_), .B1(new_n520_), .B2(KEYINPUT4), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n515_), .B1(new_n521_), .B2(new_n514_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G29gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT99), .B(G85gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT0), .B(G57gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR4_X1   g330(.A1(new_n427_), .A2(new_n454_), .A3(new_n509_), .A4(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n509_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n395_), .B(new_n534_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n531_), .B(new_n535_), .C1(new_n416_), .C2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n521_), .A2(new_n514_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n527_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT100), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT100), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n527_), .B(new_n540_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n511_), .A2(KEYINPUT4), .A3(new_n512_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n519_), .A2(new_n516_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n514_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n513_), .A2(new_n514_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n543_), .B(new_n528_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n542_), .B1(new_n544_), .B2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n536_), .B1(new_n552_), .B2(KEYINPUT101), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT101), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n554_), .B(new_n551_), .C1(new_n424_), .C2(new_n422_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n533_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT103), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n533_), .B(KEYINPUT103), .C1(new_n553_), .C2(new_n555_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n531_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n426_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n454_), .A2(KEYINPUT84), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n454_), .A2(KEYINPUT84), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n532_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n231_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n568_), .A2(new_n268_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n268_), .A2(new_n230_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n268_), .B(new_n230_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G113gat), .B(G141gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT76), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G169gat), .B(G197gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n575_), .B2(new_n572_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT77), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(KEYINPUT77), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n567_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n317_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n531_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n590_), .A2(G1gat), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n260_), .A2(KEYINPUT105), .A3(new_n250_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT105), .B1(new_n260_), .B2(new_n250_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n567_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n598_), .A2(new_n587_), .A3(new_n315_), .A4(new_n293_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G1gat), .B1(new_n599_), .B2(new_n591_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n593_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n600_), .A3(new_n601_), .ZN(G1324gat));
  OAI21_X1  g401(.A(G8gat), .B1(new_n599_), .B2(new_n426_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT39), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n590_), .A2(G8gat), .A3(new_n426_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g406(.A1(new_n590_), .A2(G15gat), .A3(new_n566_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT106), .ZN(new_n609_));
  OAI21_X1  g408(.A(G15gat), .B1(new_n599_), .B2(new_n566_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT41), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(KEYINPUT41), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n611_), .A3(new_n612_), .ZN(G1326gat));
  OAI21_X1  g412(.A(G22gat), .B1(new_n599_), .B2(new_n533_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n533_), .A2(G22gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n590_), .B2(new_n616_), .ZN(G1327gat));
  OAI21_X1  g416(.A(KEYINPUT43), .B1(new_n567_), .B2(new_n262_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT43), .ZN(new_n619_));
  INV_X1    g418(.A(new_n262_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n556_), .A2(new_n557_), .B1(new_n560_), .B2(new_n426_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n565_), .B1(new_n621_), .B2(new_n559_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n619_), .B(new_n620_), .C1(new_n622_), .C2(new_n532_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n315_), .A2(new_n587_), .A3(new_n292_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT107), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT44), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n625_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT107), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n629_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(KEYINPUT44), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(G29gat), .A3(new_n531_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n589_), .A2(new_n315_), .A3(new_n292_), .A4(new_n597_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n591_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(G1328gat));
  NOR3_X1   g439(.A1(new_n638_), .A2(G36gat), .A3(new_n426_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT45), .Z(new_n642_));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n426_), .B1(new_n630_), .B2(KEYINPUT44), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n633_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT107), .B(new_n625_), .C1(new_n618_), .C2(new_n623_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n643_), .B(new_n644_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G36gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n642_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n642_), .B(KEYINPUT46), .C1(new_n645_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NOR3_X1   g453(.A1(new_n638_), .A2(G43gat), .A3(new_n566_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n454_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n633_), .A2(new_n656_), .A3(new_n634_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n657_), .B2(G43gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n655_), .B(new_n661_), .C1(new_n657_), .C2(G43gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1330gat));
  NAND3_X1  g462(.A1(new_n635_), .A2(G50gat), .A3(new_n509_), .ZN(new_n664_));
  INV_X1    g463(.A(G50gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n638_), .B2(new_n533_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1331gat));
  NOR2_X1   g466(.A1(new_n567_), .A2(new_n587_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT110), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(KEYINPUT110), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n315_), .A3(new_n295_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n531_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n587_), .A2(new_n292_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n598_), .A2(new_n316_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G57gat), .B1(new_n676_), .B2(new_n591_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(G1332gat));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n672_), .A2(new_n679_), .A3(new_n427_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G64gat), .B1(new_n676_), .B2(new_n426_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT48), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1333gat));
  INV_X1    g482(.A(G71gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n684_), .A3(new_n565_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G71gat), .B1(new_n676_), .B2(new_n566_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT49), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1334gat));
  INV_X1    g487(.A(G78gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n672_), .A2(new_n689_), .A3(new_n509_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G78gat), .B1(new_n676_), .B2(new_n533_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT50), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1335gat));
  NOR3_X1   g492(.A1(new_n315_), .A2(new_n587_), .A3(new_n293_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n618_), .A2(new_n623_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT111), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT111), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G85gat), .B1(new_n698_), .B2(new_n591_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n597_), .ZN(new_n700_));
  NOR4_X1   g499(.A1(new_n671_), .A2(new_n315_), .A3(new_n293_), .A4(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n210_), .A3(new_n531_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(G1336gat));
  OAI21_X1  g502(.A(G92gat), .B1(new_n698_), .B2(new_n426_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n701_), .A2(new_n211_), .A3(new_n427_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1337gat));
  INV_X1    g505(.A(KEYINPUT51), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT112), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n656_), .A2(new_n205_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n701_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G99gat), .B1(new_n698_), .B2(new_n566_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(KEYINPUT112), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1338gat));
  NAND3_X1  g514(.A1(new_n701_), .A2(new_n206_), .A3(new_n509_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n694_), .A2(new_n509_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT113), .B1(new_n695_), .B2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n206_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n718_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n716_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT53), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n716_), .B(new_n727_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1339gat));
  INV_X1    g528(.A(KEYINPUT120), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n533_), .A2(new_n426_), .A3(new_n656_), .A4(new_n531_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT118), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n303_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n301_), .A2(new_n302_), .A3(new_n297_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n309_), .B1(new_n303_), .B2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n738_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(KEYINPUT116), .A3(new_n740_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n585_), .A2(new_n586_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n580_), .B1(new_n573_), .B2(new_n571_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n569_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n310_), .A2(new_n581_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n700_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT117), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n597_), .B1(new_n747_), .B2(new_n751_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT117), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n741_), .A2(new_n743_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n581_), .A2(new_n750_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT58), .B1(new_n760_), .B2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n262_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(KEYINPUT58), .A3(new_n762_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n753_), .A2(new_n754_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n293_), .B1(new_n759_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n675_), .B(KEYINPUT114), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n315_), .A3(new_n262_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n770_));
  XOR2_X1   g569(.A(new_n769_), .B(new_n770_), .Z(new_n771_));
  OAI211_X1 g570(.A(new_n732_), .B(new_n733_), .C1(new_n767_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n732_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n758_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n757_), .B1(new_n756_), .B2(KEYINPUT57), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n766_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n292_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n769_), .B(new_n770_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n773_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT59), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n772_), .B(new_n587_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G113gat), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n587_), .A2(new_n444_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n773_), .B(new_n784_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n730_), .B1(new_n783_), .B2(new_n786_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT120), .B(new_n785_), .C1(new_n782_), .C2(G113gat), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1340gat));
  OAI21_X1  g588(.A(new_n442_), .B1(new_n315_), .B2(KEYINPUT60), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n779_), .B(new_n790_), .C1(KEYINPUT60), .C2(new_n442_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT121), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n772_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G120gat), .B1(new_n793_), .B2(new_n315_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1341gat));
  OAI21_X1  g594(.A(G127gat), .B1(new_n793_), .B2(new_n292_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n439_), .A3(new_n293_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1342gat));
  OAI21_X1  g597(.A(G134gat), .B1(new_n793_), .B2(new_n262_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n779_), .A2(new_n437_), .A3(new_n597_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1343gat));
  NAND2_X1  g600(.A1(new_n777_), .A2(new_n778_), .ZN(new_n802_));
  NOR4_X1   g601(.A1(new_n565_), .A2(new_n533_), .A3(new_n591_), .A4(new_n427_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n588_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(new_n456_), .ZN(G1344gat));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n315_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(new_n457_), .ZN(G1345gat));
  OAI21_X1  g607(.A(KEYINPUT122), .B1(new_n804_), .B2(new_n292_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n802_), .A2(new_n810_), .A3(new_n293_), .A4(new_n803_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT61), .B(G155gat), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1346gat));
  OAI21_X1  g613(.A(G162gat), .B1(new_n804_), .B2(new_n262_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n597_), .A2(new_n470_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n804_), .B2(new_n816_), .ZN(G1347gat));
  NAND3_X1  g616(.A1(new_n565_), .A2(new_n591_), .A3(new_n427_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT123), .Z(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n509_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n802_), .A2(new_n587_), .A3(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT62), .B1(new_n821_), .B2(KEYINPUT22), .ZN(new_n822_));
  OAI21_X1  g621(.A(G169gat), .B1(new_n821_), .B2(KEYINPUT62), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n358_), .B2(new_n822_), .ZN(G1348gat));
  NAND2_X1  g624(.A1(new_n802_), .A2(new_n820_), .ZN(new_n826_));
  OAI22_X1  g625(.A1(new_n826_), .A2(new_n315_), .B1(KEYINPUT124), .B2(new_n359_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n359_), .A2(KEYINPUT124), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT125), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n827_), .B(new_n829_), .ZN(G1349gat));
  NOR2_X1   g629(.A1(new_n826_), .A2(new_n292_), .ZN(new_n831_));
  MUX2_X1   g630(.A(G183gat), .B(new_n384_), .S(new_n831_), .Z(G1350gat));
  OAI21_X1  g631(.A(G190gat), .B1(new_n826_), .B2(new_n262_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n597_), .A2(new_n385_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT126), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n826_), .B2(new_n835_), .ZN(G1351gat));
  NOR4_X1   g635(.A1(new_n565_), .A2(new_n533_), .A3(new_n531_), .A4(new_n426_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n802_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n588_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n323_), .ZN(G1352gat));
  NOR2_X1   g639(.A1(new_n838_), .A2(new_n315_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(G204gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n319_), .A2(new_n321_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n841_), .ZN(G1353gat));
  AOI21_X1  g643(.A(new_n292_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n802_), .A2(new_n837_), .A3(new_n845_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n846_), .A2(KEYINPUT127), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(KEYINPUT127), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n850_));
  INV_X1    g649(.A(G211gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n847_), .A2(new_n850_), .A3(new_n851_), .A4(new_n848_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1354gat));
  OAI21_X1  g654(.A(G218gat), .B1(new_n838_), .B2(new_n262_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n700_), .A2(G218gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n838_), .B2(new_n857_), .ZN(G1355gat));
endmodule


