//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .A4(KEYINPUT87), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  OAI22_X1  g006(.A1(new_n207_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n206_), .A2(new_n208_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n221_), .A2(KEYINPUT88), .A3(new_n208_), .A4(new_n206_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n216_), .A2(KEYINPUT1), .B1(new_n204_), .B2(new_n205_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n209_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT83), .B(G127gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G113gat), .ZN(new_n231_));
  INV_X1    g030(.A(G120gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G134gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n230_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n238_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n229_), .A3(new_n236_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n228_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n223_), .A3(new_n227_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT4), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n228_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT97), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(new_n245_), .A3(new_n249_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT97), .A4(new_n250_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G1gat), .B(G29gat), .ZN(new_n257_));
  INV_X1    g056(.A(G85gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G57gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .A4(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT78), .B(G183gat), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(KEYINPUT25), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT26), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT79), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT79), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT26), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n274_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n273_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT79), .B(KEYINPUT26), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n273_), .A2(new_n274_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n272_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT24), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n269_), .B1(new_n285_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT82), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n291_), .B1(new_n296_), .B2(KEYINPUT23), .ZN(new_n297_));
  NOR3_X1   g096(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n289_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n280_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(new_n282_), .B2(new_n274_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n302_), .A2(new_n273_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n303_));
  OAI211_X1 g102(.A(KEYINPUT81), .B(new_n300_), .C1(new_n303_), .C2(new_n272_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n290_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT30), .ZN(new_n306_));
  INV_X1    g105(.A(new_n286_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT22), .B(G169gat), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n293_), .A2(new_n295_), .A3(KEYINPUT23), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n292_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n271_), .A2(G190gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n310_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n305_), .A2(new_n306_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n306_), .B1(new_n305_), .B2(new_n316_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G15gat), .B(G43gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(G71gat), .B(G99gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n317_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n305_), .A2(new_n316_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT30), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n305_), .A2(new_n306_), .A3(new_n316_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n323_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n268_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n324_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT85), .A3(new_n268_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n334_), .A3(new_n267_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT84), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT84), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n333_), .A2(new_n334_), .A3(new_n340_), .A4(new_n267_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n337_), .A2(KEYINPUT86), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT86), .B1(new_n337_), .B2(new_n342_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n266_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT93), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT90), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n352_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n351_), .A2(new_n355_), .A3(new_n352_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(KEYINPUT92), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n350_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n350_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n228_), .B2(KEYINPUT29), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n358_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT91), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(KEYINPUT91), .A3(new_n358_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n348_), .B1(new_n371_), .B2(KEYINPUT94), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n362_), .A2(new_n363_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n365_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n366_), .A2(KEYINPUT91), .A3(new_n358_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT91), .B1(new_n366_), .B2(new_n358_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT89), .B1(new_n377_), .B2(new_n347_), .ZN(new_n378_));
  OR3_X1    g177(.A1(new_n228_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT28), .B(G22gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(G50gat), .B1(new_n228_), .B2(KEYINPUT29), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n381_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n372_), .A2(new_n378_), .A3(new_n382_), .A4(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n382_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n371_), .A2(new_n348_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(KEYINPUT89), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n348_), .B(new_n371_), .C1(new_n387_), .C2(KEYINPUT94), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n286_), .A2(KEYINPUT95), .A3(KEYINPUT24), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT95), .B1(new_n286_), .B2(KEYINPUT24), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n288_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(new_n314_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT26), .B(G190gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n298_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n291_), .B(new_n401_), .C1(new_n296_), .C2(KEYINPUT23), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n397_), .A2(new_n400_), .B1(new_n402_), .B2(new_n310_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n356_), .A2(new_n357_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n393_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n310_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n395_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n288_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n286_), .A2(KEYINPUT95), .A3(KEYINPUT24), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(new_n400_), .A3(new_n313_), .A4(new_n311_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(KEYINPUT96), .A3(new_n358_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n392_), .B1(new_n405_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n305_), .A2(new_n316_), .A3(new_n404_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT19), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G92gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT18), .B(G64gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n326_), .A2(new_n358_), .ZN(new_n424_));
  AOI211_X1 g223(.A(new_n392_), .B(new_n418_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n423_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n418_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n425_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n404_), .B1(new_n305_), .B2(new_n316_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n428_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT100), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n412_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n418_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n414_), .A2(new_n415_), .A3(new_n429_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n428_), .ZN(new_n443_));
  AND4_X1   g242(.A1(new_n438_), .A2(new_n443_), .A3(KEYINPUT27), .A4(new_n427_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n416_), .A2(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n423_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n438_), .B1(new_n447_), .B2(new_n443_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n391_), .B(new_n437_), .C1(new_n444_), .C2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n202_), .B1(new_n345_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT85), .B1(new_n335_), .B2(new_n268_), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n331_), .B(new_n267_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n339_), .A2(new_n341_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n337_), .A2(KEYINPUT86), .A3(new_n342_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n265_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n449_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT102), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n264_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n244_), .A2(new_n464_), .A3(new_n245_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n250_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n262_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n427_), .A2(new_n434_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n461_), .B1(new_n463_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n264_), .B(KEYINPUT33), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n427_), .A2(new_n434_), .A3(new_n469_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT99), .A3(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n423_), .A2(KEYINPUT32), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n442_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n419_), .A2(new_n426_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n265_), .B(new_n476_), .C1(new_n477_), .C2(new_n475_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(new_n474_), .A3(new_n391_), .A4(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n479_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n391_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n437_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(new_n265_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n450_), .A2(new_n460_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT67), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G85gat), .B(G92gat), .Z(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT10), .B(G99gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT64), .B(G106gat), .ZN(new_n495_));
  AOI22_X1  g294(.A1(KEYINPUT9), .A2(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(KEYINPUT9), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n492_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n500_));
  NOR2_X1   g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(new_n489_), .A3(new_n491_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n493_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n507_), .A3(new_n493_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n499_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G57gat), .B(G64gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(KEYINPUT11), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G78gat), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n486_), .B1(new_n509_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT12), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G230gat), .A2(G233gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n509_), .A2(new_n516_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n492_), .A2(new_n498_), .A3(new_n496_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n504_), .A2(new_n507_), .A3(new_n493_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n507_), .B1(new_n504_), .B2(new_n493_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT12), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n486_), .A3(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n520_), .A2(new_n526_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n519_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n485_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n485_), .B2(new_n532_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT69), .B(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT5), .B(G176gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G120gat), .B(G148gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n537_), .B(new_n538_), .Z(new_n539_));
  OR2_X1    g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(new_n539_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n541_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(KEYINPUT13), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G29gat), .B(G36gat), .ZN(new_n550_));
  INV_X1    g349(.A(G50gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT71), .B(G43gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT15), .ZN(new_n555_));
  XOR2_X1   g354(.A(G15gat), .B(G22gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT75), .B(G1gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(G8gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n558_), .B2(KEYINPUT14), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G1gat), .B(G8gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n554_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n561_), .B(new_n554_), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(G229gat), .A3(G233gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n484_), .A2(new_n549_), .A3(new_n578_), .ZN(new_n579_));
  MUX2_X1   g378(.A(new_n554_), .B(new_n555_), .S(new_n524_), .Z(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n580_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(KEYINPUT35), .A3(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT74), .ZN(new_n588_));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT36), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n585_), .A2(new_n593_), .A3(new_n586_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT72), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n585_), .A2(new_n586_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT73), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n587_), .A2(new_n592_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n604_), .B(new_n605_), .C1(new_n603_), .C2(new_n599_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n516_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n563_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n610_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n610_), .A2(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT77), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT77), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n607_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n579_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n557_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n265_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT38), .ZN(new_n630_));
  INV_X1    g429(.A(new_n600_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(new_n625_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n579_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n634_), .B2(new_n266_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n630_), .A2(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(G8gat), .ZN(new_n637_));
  AND2_X1   g436(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n638_));
  AOI211_X1 g437(.A(new_n637_), .B(new_n638_), .C1(new_n633_), .C2(new_n482_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n627_), .A2(new_n637_), .A3(new_n482_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n456_), .A2(new_n457_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n633_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n627_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n633_), .B2(new_n481_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n627_), .A2(new_n652_), .A3(new_n481_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(new_n607_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n484_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n646_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n483_), .A3(new_n479_), .ZN(new_n661_));
  AND4_X1   g460(.A1(KEYINPUT102), .A2(new_n646_), .A3(new_n266_), .A4(new_n459_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n458_), .B2(new_n459_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT43), .B1(new_n664_), .B2(new_n607_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n659_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n549_), .A2(new_n578_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n667_), .A4(new_n625_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n657_), .B1(new_n484_), .B2(new_n658_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(KEYINPUT43), .A3(new_n607_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n667_), .A4(new_n625_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n668_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n266_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n631_), .A2(new_n625_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT105), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n579_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT106), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n266_), .A2(G29gat), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n682_), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n668_), .A2(new_n482_), .A3(new_n673_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT108), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n668_), .A2(new_n686_), .A3(new_n482_), .A4(new_n673_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(G36gat), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n685_), .A2(new_n690_), .A3(G36gat), .A4(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n482_), .B(KEYINPUT110), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n679_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n679_), .A2(new_n697_), .A3(new_n693_), .A4(new_n694_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n696_), .A2(new_n698_), .B1(KEYINPUT111), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n692_), .A2(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n699_), .A2(KEYINPUT111), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT112), .Z(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n692_), .A2(new_n703_), .A3(new_n700_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n674_), .B2(new_n660_), .ZN(new_n708_));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n679_), .A2(new_n709_), .A3(new_n646_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g511(.A(G50gat), .B1(new_n674_), .B2(new_n391_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n679_), .A2(new_n551_), .A3(new_n481_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1331gat));
  NOR3_X1   g514(.A1(new_n484_), .A2(new_n577_), .A3(new_n548_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n632_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n266_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n626_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT113), .Z(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n265_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n719_), .B1(new_n722_), .B2(new_n718_), .ZN(G1332gat));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(new_n724_), .A3(new_n694_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n694_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G64gat), .B1(new_n717_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT48), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT114), .Z(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n721_), .A2(new_n731_), .A3(new_n646_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G71gat), .B1(new_n717_), .B2(new_n660_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT49), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1334gat));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n721_), .A2(new_n736_), .A3(new_n481_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G78gat), .B1(new_n717_), .B2(new_n391_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT115), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT115), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n739_), .A2(new_n740_), .A3(KEYINPUT50), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n737_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT116), .Z(G1335gat));
  NAND2_X1  g545(.A1(new_n716_), .A2(new_n677_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n265_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n625_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n659_), .A2(new_n665_), .A3(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n548_), .A2(new_n577_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n266_), .A2(new_n258_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n749_), .B1(new_n754_), .B2(new_n755_), .ZN(G1336gat));
  AOI21_X1  g555(.A(G92gat), .B1(new_n748_), .B2(new_n482_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n694_), .A2(G92gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n754_), .B2(new_n758_), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n753_), .B2(new_n660_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n748_), .A2(new_n494_), .A3(new_n646_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g562(.A(G106gat), .B1(new_n753_), .B2(new_n391_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT52), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(KEYINPUT52), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n481_), .A2(new_n495_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n765_), .A2(new_n766_), .B1(new_n748_), .B2(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n768_), .B(new_n769_), .Z(G1339gat));
  NOR3_X1   g569(.A1(new_n660_), .A2(new_n266_), .A3(new_n449_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT120), .ZN(new_n772_));
  INV_X1    g571(.A(new_n539_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n518_), .A2(new_n520_), .A3(new_n528_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n531_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n529_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n775_), .A2(new_n774_), .A3(new_n531_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT56), .B(new_n773_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n527_), .B1(new_n526_), .B2(new_n486_), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n524_), .C2(new_n525_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n519_), .B1(new_n785_), .B2(new_n520_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n529_), .B1(new_n786_), .B2(new_n774_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n779_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n789_), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(new_n773_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n773_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n782_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n541_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n578_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n568_), .A2(new_n566_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n565_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n573_), .B(new_n800_), .C1(new_n801_), .C2(new_n566_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n576_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n545_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n794_), .A2(new_n796_), .A3(KEYINPUT119), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n799_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n600_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n772_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT120), .B(KEYINPUT57), .C1(new_n807_), .C2(new_n600_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n773_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n795_), .B1(new_n813_), .B2(KEYINPUT121), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n793_), .A2(new_n815_), .A3(new_n780_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n804_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n816_), .A4(new_n804_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n607_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT122), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n819_), .A2(new_n607_), .A3(new_n820_), .A4(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n794_), .A2(new_n796_), .A3(KEYINPUT119), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT119), .B1(new_n794_), .B2(new_n796_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n631_), .B1(new_n827_), .B2(new_n805_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n822_), .A2(new_n824_), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n750_), .B1(new_n812_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n626_), .A2(new_n548_), .A3(new_n578_), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT54), .Z(new_n832_));
  OAI21_X1  g631(.A(new_n771_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834_), .B2(new_n577_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n832_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT123), .B(new_n821_), .C1(new_n828_), .C2(KEYINPUT57), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n807_), .B2(new_n600_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n821_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n828_), .A2(KEYINPUT57), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n837_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n836_), .B1(new_n843_), .B2(new_n750_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n660_), .A2(KEYINPUT59), .A3(new_n266_), .A4(new_n449_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n833_), .A2(KEYINPUT59), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n578_), .A2(new_n231_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n835_), .B1(new_n846_), .B2(new_n847_), .ZN(G1340gat));
  OAI21_X1  g647(.A(new_n232_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n834_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n232_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n846_), .A2(new_n549_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n232_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n834_), .B2(new_n750_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n750_), .A2(G127gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n846_), .B2(new_n854_), .ZN(G1342gat));
  AOI21_X1  g654(.A(new_n234_), .B1(new_n846_), .B2(new_n607_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n833_), .A2(G134gat), .A3(new_n600_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT124), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n844_), .A2(new_n845_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n607_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G134gat), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(new_n857_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n858_), .A2(new_n865_), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n812_), .A2(new_n829_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n832_), .B1(new_n867_), .B2(new_n625_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n646_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n869_), .A2(new_n265_), .A3(new_n481_), .A4(new_n726_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n204_), .A3(new_n577_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G141gat), .B1(new_n870_), .B2(new_n578_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1344gat));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n205_), .A3(new_n549_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G148gat), .B1(new_n870_), .B2(new_n548_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1345gat));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n871_), .B2(new_n750_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n878_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n870_), .A2(new_n625_), .A3(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n870_), .A2(new_n883_), .A3(new_n658_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n871_), .A2(new_n631_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(G1347gat));
  NOR3_X1   g685(.A1(new_n726_), .A2(new_n265_), .A3(new_n660_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n844_), .A2(new_n391_), .A3(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888_), .B2(new_n578_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n308_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n888_), .A2(new_n578_), .A3(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT62), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1348gat));
  INV_X1    g695(.A(new_n888_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G176gat), .B1(new_n897_), .B2(new_n549_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n868_), .A2(new_n481_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n899_), .A2(G176gat), .A3(new_n887_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n549_), .B2(new_n900_), .ZN(G1349gat));
  INV_X1    g700(.A(new_n398_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n902_), .A3(new_n750_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT125), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n897_), .A2(new_n905_), .A3(new_n902_), .A4(new_n750_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n899_), .A2(new_n750_), .A3(new_n887_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n271_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n904_), .A2(new_n906_), .A3(new_n909_), .ZN(G1350gat));
  NAND3_X1  g709(.A1(new_n897_), .A2(new_n399_), .A3(new_n631_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G190gat), .B1(new_n888_), .B2(new_n658_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1351gat));
  NOR2_X1   g712(.A1(new_n726_), .A2(new_n265_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n869_), .A2(new_n481_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n577_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G197gat), .ZN(new_n917_));
  INV_X1    g716(.A(G197gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n915_), .A2(new_n918_), .A3(new_n577_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1352gat));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(G204gat), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(G204gat), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n915_), .B(new_n549_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n915_), .A2(new_n549_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n922_), .ZN(G1353gat));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927_));
  INV_X1    g726(.A(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n625_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n915_), .A2(new_n929_), .A3(new_n933_), .A4(new_n934_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n869_), .A2(new_n481_), .A3(new_n914_), .A4(new_n934_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n927_), .B(new_n928_), .C1(new_n936_), .C2(new_n932_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1354gat));
  NAND2_X1  g737(.A1(new_n915_), .A2(new_n631_), .ZN(new_n939_));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n658_), .A2(new_n940_), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n939_), .A2(new_n940_), .B1(new_n915_), .B2(new_n941_), .ZN(G1355gat));
endmodule


