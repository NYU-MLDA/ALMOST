//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(new_n203_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT87), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n202_), .A2(new_n203_), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n205_), .B(new_n204_), .C1(new_n210_), .C2(KEYINPUT87), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(KEYINPUT26), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT77), .A3(G190gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G169gat), .ZN(new_n226_));
  INV_X1    g025(.A(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT24), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n220_), .A2(new_n225_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT78), .B(new_n230_), .C1(new_n235_), .C2(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  AOI21_X1  g036(.A(G176gat), .B1(new_n233_), .B2(new_n234_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n230_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n223_), .B(new_n224_), .C1(G183gat), .C2(G190gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n212_), .A2(new_n232_), .A3(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n241_), .B(new_n230_), .C1(new_n235_), .C2(G176gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT26), .B(G190gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n213_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n211_), .A3(new_n209_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n250_), .A3(KEYINPUT20), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n209_), .A2(new_n211_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n242_), .A2(new_n232_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n245_), .A2(new_n248_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n212_), .A2(new_n244_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n253_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n257_), .A2(KEYINPUT20), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G64gat), .B(G92gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n254_), .A2(new_n269_), .A3(new_n261_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT27), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n243_), .A2(KEYINPUT20), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(KEYINPUT94), .A3(new_n260_), .A4(new_n250_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n257_), .A2(KEYINPUT20), .A3(new_n259_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(new_n253_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n251_), .A2(new_n253_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n274_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n267_), .B(KEYINPUT97), .Z(new_n280_));
  AOI21_X1  g079(.A(new_n272_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n271_), .B1(new_n281_), .B2(KEYINPUT27), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G228gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n285_));
  INV_X1    g084(.A(G141gat), .ZN(new_n286_));
  INV_X1    g085(.A(G148gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT3), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(G141gat), .B2(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT83), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(KEYINPUT83), .A3(new_n293_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT2), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n291_), .A2(new_n296_), .A3(new_n297_), .A4(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT81), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G155gat), .A3(G162gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT84), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n303_), .A2(new_n305_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT82), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n301_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n303_), .A2(new_n305_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(KEYINPUT1), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n298_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n285_), .B1(new_n311_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n284_), .B1(new_n323_), .B2(new_n212_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n300_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n309_), .B1(new_n300_), .B2(new_n306_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n321_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n317_), .B1(new_n316_), .B2(KEYINPUT1), .ZN(new_n329_));
  AOI211_X1 g128(.A(KEYINPUT82), .B(new_n313_), .C1(new_n303_), .C2(new_n305_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n328_), .B1(new_n331_), .B2(new_n315_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT29), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n283_), .A3(new_n255_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n324_), .A2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G78gat), .B(G106gat), .Z(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(KEYINPUT89), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n337_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G22gat), .B(G50gat), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n311_), .A2(new_n322_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(KEYINPUT29), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n343_));
  INV_X1    g142(.A(new_n340_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n311_), .A2(new_n322_), .A3(new_n285_), .A4(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n343_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n338_), .B(new_n339_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n335_), .A2(KEYINPUT88), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n324_), .A2(new_n334_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n336_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT86), .B1(new_n347_), .B2(new_n348_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n348_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n346_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n335_), .A2(KEYINPUT88), .A3(new_n336_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n354_), .A2(new_n355_), .A3(new_n358_), .A4(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n282_), .A2(new_n349_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT99), .ZN(new_n362_));
  XOR2_X1   g161(.A(G127gat), .B(G134gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G113gat), .B(G120gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n365_), .A2(new_n368_), .A3(KEYINPUT80), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT80), .B1(new_n365_), .B2(new_n368_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n365_), .A2(new_n368_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n311_), .A2(new_n322_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n372_), .A2(new_n377_), .A3(new_n378_), .A4(KEYINPUT4), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n372_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT92), .B1(new_n372_), .B2(KEYINPUT4), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n372_), .A2(new_n377_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n384_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n369_), .A2(new_n370_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n311_), .B2(new_n322_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n372_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n383_), .B1(new_n400_), .B2(new_n379_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n394_), .B1(new_n401_), .B2(new_n387_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT95), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n393_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n385_), .A2(KEYINPUT95), .A3(new_n388_), .A4(new_n392_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n371_), .B(KEYINPUT31), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n256_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n411_));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G71gat), .B(G99gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n410_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT99), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n282_), .A2(new_n360_), .A3(new_n417_), .A4(new_n349_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n362_), .A2(new_n406_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT100), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n360_), .A2(new_n349_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n406_), .A2(new_n421_), .A3(new_n282_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT98), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT96), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n279_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n262_), .A2(new_n426_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n404_), .A2(new_n405_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n386_), .A2(new_n383_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n384_), .B1(new_n400_), .B2(new_n379_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n382_), .A2(new_n383_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT93), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n435_), .A3(new_n394_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n393_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n268_), .A2(new_n270_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n385_), .A2(KEYINPUT33), .A3(new_n388_), .A4(new_n392_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n429_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n421_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n425_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI211_X1 g244(.A(KEYINPUT96), .B(new_n421_), .C1(new_n429_), .C2(new_n441_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n424_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n416_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n420_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G43gat), .B(G50gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n454_), .B1(new_n465_), .B2(KEYINPUT74), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n461_), .A2(new_n464_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(KEYINPUT74), .A3(new_n454_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n453_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n464_), .B(KEYINPUT15), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n461_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n465_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n452_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G169gat), .B(G197gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n474_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n474_), .B2(new_n480_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n451_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n474_), .A2(new_n480_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n483_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n485_), .A3(KEYINPUT76), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G71gat), .B(G78gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(KEYINPUT11), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n498_), .B2(new_n495_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT10), .B(G99gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT64), .ZN(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT9), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G85gat), .A3(G92gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n507_));
  AND2_X1   g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G85gat), .B(G92gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n504_), .A2(new_n506_), .A3(new_n509_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n508_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n515_), .B(KEYINPUT67), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n508_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT7), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n514_), .B1(new_n524_), .B2(new_n511_), .ZN(new_n525_));
  AOI211_X1 g324(.A(KEYINPUT8), .B(new_n510_), .C1(new_n509_), .C2(new_n523_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n513_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT68), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n529_), .B(new_n513_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n500_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT12), .B1(new_n527_), .B2(new_n499_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n499_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n527_), .B(new_n499_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G176gat), .B(G204gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(new_n540_), .A3(new_n546_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n541_), .A2(KEYINPUT70), .A3(new_n547_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n551_), .A2(new_n552_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n556_), .A3(new_n552_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n492_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n450_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n475_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT35), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n527_), .A2(new_n464_), .B1(KEYINPUT35), .B2(new_n565_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n563_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT36), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n571_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n574_), .B(KEYINPUT36), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n562_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n577_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n584_), .B2(new_n570_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n578_), .A3(new_n561_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n461_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n500_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  XOR2_X1   g391(.A(G183gat), .B(G211gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n592_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n587_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n560_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n406_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n456_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT38), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n579_), .A2(new_n582_), .A3(KEYINPUT101), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT101), .B1(new_n579_), .B2(new_n582_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n602_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n560_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(new_n605_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n456_), .B2(new_n614_), .ZN(G1324gat));
  INV_X1    g414(.A(new_n282_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n457_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT39), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n604_), .A2(new_n457_), .A3(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n613_), .B2(new_n416_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT41), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n604_), .A2(new_n622_), .A3(new_n416_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  INV_X1    g425(.A(G22gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n613_), .B2(new_n421_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT42), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n604_), .A2(new_n627_), .A3(new_n421_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1327gat));
  NOR2_X1   g430(.A1(new_n610_), .A2(new_n601_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n444_), .A2(new_n446_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n416_), .B1(new_n633_), .B2(new_n424_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n558_), .B(new_n632_), .C1(new_n634_), .C2(new_n420_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT102), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n419_), .B(KEYINPUT100), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n422_), .B(KEYINPUT98), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n639_), .B2(new_n416_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n558_), .A4(new_n632_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(G29gat), .B1(new_n644_), .B2(new_n605_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n558_), .A2(new_n602_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n587_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT43), .B1(new_n450_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n649_), .B(new_n587_), .C1(new_n634_), .C2(new_n420_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n646_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(G29gat), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n653_), .B(new_n646_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n406_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n645_), .B1(new_n655_), .B2(new_n657_), .ZN(G1328gat));
  NOR2_X1   g457(.A1(new_n282_), .A2(G36gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n636_), .A2(new_n642_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n636_), .A2(new_n642_), .A3(new_n662_), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n616_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n667_));
  OAI21_X1  g466(.A(G36gat), .B1(new_n667_), .B2(new_n656_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(KEYINPUT45), .A3(new_n663_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n666_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT104), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n666_), .A2(new_n668_), .A3(new_n673_), .A4(new_n669_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n670_), .A2(new_n672_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n671_), .A2(new_n678_), .A3(new_n672_), .A4(new_n674_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n677_), .A3(new_n679_), .ZN(G1329gat));
  NAND2_X1  g479(.A1(new_n654_), .A2(G43gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n416_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n643_), .A2(new_n449_), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n681_), .A2(new_n682_), .B1(G43gat), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n644_), .B2(new_n421_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n654_), .A2(G50gat), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n656_), .A2(new_n443_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n687_), .B2(new_n688_), .ZN(G1331gat));
  INV_X1    g488(.A(new_n492_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n554_), .A2(new_n557_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n450_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(new_n603_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n605_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n692_), .A2(new_n612_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(G57gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n605_), .B2(new_n696_), .ZN(G1332gat));
  INV_X1    g496(.A(G64gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n695_), .B2(new_n616_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT48), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(new_n698_), .A3(new_n616_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n695_), .B2(new_n416_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT106), .Z(new_n705_));
  INV_X1    g504(.A(KEYINPUT49), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n693_), .A2(new_n416_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n707_), .B(new_n708_), .C1(G71gat), .C2(new_n709_), .ZN(G1334gat));
  INV_X1    g509(.A(G78gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n695_), .B2(new_n421_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT50), .Z(new_n713_));
  NAND2_X1  g512(.A1(new_n421_), .A2(new_n711_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n693_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1335gat));
  AND2_X1   g516(.A1(new_n692_), .A2(new_n632_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n605_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n691_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n602_), .A3(new_n492_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT108), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n648_), .A2(new_n650_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT109), .Z(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(G85gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n719_), .B1(new_n726_), .B2(new_n605_), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n718_), .B2(new_n616_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n725_), .A2(new_n616_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n416_), .A3(new_n723_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n416_), .A2(new_n502_), .ZN(new_n732_));
  AOI22_X1  g531(.A1(new_n731_), .A2(G99gat), .B1(new_n718_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(G1338gat));
  NAND3_X1  g534(.A1(new_n722_), .A2(new_n421_), .A3(new_n723_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G106gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(KEYINPUT111), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT111), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n738_), .A2(KEYINPUT111), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n736_), .A2(G106gat), .A3(new_n740_), .A4(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n718_), .A2(new_n503_), .A3(new_n421_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(G1339gat));
  AND3_X1   g545(.A1(new_n362_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n488_), .A2(new_n491_), .A3(new_n601_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n583_), .A2(new_n586_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n749_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n557_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n750_), .B(new_n752_), .C1(new_n753_), .C2(new_n553_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT115), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n754_), .A2(KEYINPUT114), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n760_), .A3(new_n756_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n759_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n759_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT115), .B(KEYINPUT54), .C1(new_n754_), .C2(KEYINPUT114), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n762_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT55), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n532_), .A2(new_n533_), .A3(new_n536_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n531_), .A2(KEYINPUT12), .B1(new_n535_), .B2(new_n534_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n533_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT12), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n776_), .B(new_n500_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n536_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT116), .B(new_n539_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n774_), .A2(new_n768_), .A3(KEYINPUT55), .A4(new_n533_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n772_), .A2(new_n775_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n547_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n492_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n786_), .A4(new_n547_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n784_), .A2(new_n550_), .A3(new_n785_), .A4(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n473_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n453_), .B1(new_n789_), .B2(new_n471_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n483_), .B1(new_n478_), .B2(new_n452_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT119), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n452_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  INV_X1    g593(.A(new_n791_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n485_), .A3(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT120), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n788_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT57), .B1(new_n800_), .B2(new_n610_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n802_), .B(new_n611_), .C1(new_n788_), .C2(new_n799_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n781_), .A2(new_n786_), .A3(new_n547_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n785_), .A2(new_n550_), .A3(new_n798_), .A4(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n805_), .A2(new_n550_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(KEYINPUT58), .A3(new_n798_), .A4(new_n785_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n808_), .A2(new_n810_), .A3(new_n587_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n601_), .B1(new_n804_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n605_), .B(new_n747_), .C1(new_n767_), .C2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815_), .B2(new_n690_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(KEYINPUT59), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n801_), .A2(new_n803_), .A3(new_n811_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n762_), .B(new_n766_), .C1(new_n818_), .C2(new_n601_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n605_), .A4(new_n747_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n822_), .A2(new_n690_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n823_), .B2(G113gat), .ZN(G1340gat));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n720_), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G120gat), .ZN(new_n826_));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n691_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n815_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n827_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n815_), .B2(new_n601_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n601_), .A2(G127gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n822_), .B2(new_n836_), .ZN(G1342gat));
  AOI21_X1  g636(.A(G134gat), .B1(new_n815_), .B2(new_n611_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n587_), .A2(G134gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n822_), .B2(new_n839_), .ZN(G1343gat));
  AND2_X1   g639(.A1(new_n819_), .A2(new_n605_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n616_), .A2(new_n416_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n421_), .A3(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n492_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n286_), .ZN(G1344gat));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n691_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT122), .B(G148gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  INV_X1    g647(.A(new_n843_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n601_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  AOI21_X1  g651(.A(G162gat), .B1(new_n849_), .B2(new_n611_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n587_), .A2(G162gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT123), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n849_), .B2(new_n855_), .ZN(G1347gat));
  NOR2_X1   g655(.A1(new_n605_), .A2(new_n421_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n819_), .A2(new_n416_), .A3(new_n616_), .A4(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G169gat), .B1(new_n858_), .B2(new_n492_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n858_), .A2(new_n492_), .A3(new_n235_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT62), .B(G169gat), .C1(new_n858_), .C2(new_n492_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT124), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n861_), .A2(new_n866_), .A3(new_n862_), .A4(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1348gat));
  NOR2_X1   g667(.A1(new_n858_), .A2(new_n691_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n227_), .ZN(G1349gat));
  NOR2_X1   g669(.A1(new_n858_), .A2(new_n602_), .ZN(new_n871_));
  MUX2_X1   g670(.A(G183gat), .B(new_n213_), .S(new_n871_), .Z(G1350gat));
  OAI21_X1  g671(.A(G190gat), .B1(new_n858_), .B2(new_n647_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n611_), .A2(new_n246_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n858_), .B2(new_n874_), .ZN(G1351gat));
  NAND4_X1  g674(.A1(new_n819_), .A2(new_n406_), .A3(new_n421_), .A4(new_n616_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n416_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n690_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n720_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n876_), .A2(new_n416_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n602_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(KEYINPUT125), .B(new_n882_), .C1(new_n883_), .C2(new_n602_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n883_), .A2(new_n602_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT63), .B(G211gat), .Z(new_n889_));
  AOI22_X1  g688(.A1(new_n886_), .A2(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1354gat));
  NAND2_X1  g689(.A1(new_n877_), .A2(new_n611_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT126), .B(G218gat), .Z(new_n892_));
  NOR2_X1   g691(.A1(new_n647_), .A2(new_n892_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n891_), .A2(new_n892_), .B1(new_n877_), .B2(new_n893_), .ZN(G1355gat));
endmodule


