//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT85), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n212_), .A2(new_n205_), .A3(new_n204_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(new_n208_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n209_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT88), .ZN(new_n220_));
  INV_X1    g019(.A(new_n212_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(KEYINPUT88), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT87), .B(G176gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G169gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n210_), .A2(KEYINPUT86), .A3(KEYINPUT22), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n218_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT90), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  XOR2_X1   g040(.A(new_n232_), .B(new_n241_), .Z(new_n242_));
  XNOR2_X1  g041(.A(G15gat), .B(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n242_), .B(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT91), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n251_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT2), .Z(new_n256_));
  OAI21_X1  g055(.A(new_n250_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n248_), .A2(KEYINPUT1), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n259_), .A2(new_n255_), .A3(new_n251_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n239_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n235_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT4), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT101), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT101), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n263_), .A2(new_n267_), .A3(new_n264_), .A4(KEYINPUT4), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n263_), .A2(KEYINPUT4), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n263_), .A2(new_n272_), .A3(new_n264_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G57gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G85gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(G1gat), .B(G29gat), .Z(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT102), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT18), .B(G64gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(G92gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT19), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT99), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT20), .ZN(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(G197gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(KEYINPUT92), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G204gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n293_), .B1(new_n297_), .B2(G197gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT21), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n294_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT93), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n292_), .A2(G197gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT93), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n294_), .A2(new_n296_), .A3(new_n307_), .A4(new_n303_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT21), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n300_), .B1(new_n298_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(KEYINPUT94), .A3(KEYINPUT21), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT95), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n312_), .A2(new_n318_), .A3(new_n314_), .A4(new_n315_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n302_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n229_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n291_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n309_), .A2(KEYINPUT94), .A3(KEYINPUT21), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT94), .B1(new_n309_), .B2(KEYINPUT21), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n318_), .B1(new_n325_), .B2(new_n314_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n319_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n301_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n216_), .A2(new_n207_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G169gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n212_), .B1(new_n223_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n219_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n290_), .B1(new_n322_), .B2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n301_), .B(new_n333_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT20), .ZN(new_n338_));
  INV_X1    g137(.A(new_n289_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n287_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n290_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n321_), .B(new_n301_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT20), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n320_), .A2(new_n333_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n343_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n291_), .B1(new_n320_), .B2(new_n333_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n328_), .A2(new_n229_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n350_), .A3(new_n286_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(KEYINPUT100), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT100), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n287_), .C1(new_n336_), .C2(new_n341_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n282_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n270_), .A2(new_n272_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n272_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n278_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n278_), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n362_), .B(new_n357_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n349_), .B1(new_n348_), .B2(KEYINPUT103), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT103), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n338_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n289_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n345_), .A2(new_n346_), .A3(new_n343_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n286_), .A2(KEYINPUT32), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n364_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n347_), .A2(new_n350_), .A3(new_n372_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n355_), .A2(new_n361_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G78gat), .B(G106gat), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G228gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n262_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n328_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n379_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n320_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n378_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n328_), .A2(new_n379_), .A3(new_n383_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n385_), .B1(new_n320_), .B2(new_n382_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n377_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n381_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT28), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n392_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT96), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT96), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n399_), .A3(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT97), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n396_), .B1(new_n391_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n387_), .A2(KEYINPUT97), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT98), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n388_), .A2(new_n389_), .A3(new_n377_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n377_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n402_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  AND4_X1   g207(.A1(KEYINPUT98), .A2(new_n408_), .A3(new_n404_), .A4(new_n395_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n401_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT104), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n376_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n352_), .A2(new_n354_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n281_), .A3(new_n361_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n374_), .A2(new_n375_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n408_), .A2(new_n404_), .A3(new_n395_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT98), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n403_), .A2(KEYINPUT98), .A3(new_n404_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n419_), .A2(new_n420_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT104), .B1(new_n416_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n412_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n413_), .A2(KEYINPUT27), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n286_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n351_), .B1(new_n425_), .B2(KEYINPUT106), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n320_), .A2(new_n321_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n338_), .B2(new_n366_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n348_), .A2(KEYINPUT103), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n339_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(KEYINPUT106), .B(new_n287_), .C1(new_n430_), .C2(new_n369_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT27), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT107), .B1(new_n426_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n351_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n287_), .B1(new_n430_), .B2(new_n369_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT106), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT27), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n425_), .B2(KEYINPUT106), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT107), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n424_), .B1(new_n433_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT105), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n364_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n419_), .A2(new_n420_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n401_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n247_), .B1(new_n423_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n242_), .B(new_n245_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(new_n410_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n444_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n424_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n426_), .A2(new_n432_), .A3(KEYINPUT107), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n440_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT108), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n442_), .A2(KEYINPUT108), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n452_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n448_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT75), .B(G43gat), .ZN(new_n463_));
  INV_X1    g262(.A(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n466_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT81), .B(G8gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(G1gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(G1gat), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G8gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n469_), .B(KEYINPUT82), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(new_n479_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n479_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n462_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n462_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(new_n210_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(new_n303_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n492_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n495_), .B1(new_n490_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n461_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n504_), .A2(G99gat), .A3(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT7), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT6), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT8), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT10), .B(G99gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT64), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT65), .B(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT66), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n508_), .B1(KEYINPUT9), .B2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(KEYINPUT9), .B2(new_n510_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n511_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n506_), .B(KEYINPUT68), .ZN(new_n522_));
  INV_X1    g321(.A(new_n508_), .ZN(new_n523_));
  OAI211_X1 g322(.A(KEYINPUT8), .B(new_n510_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n469_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n503_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n471_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n532_), .A2(new_n533_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n527_), .A2(new_n535_), .A3(new_n536_), .A4(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT76), .B(G134gat), .ZN(new_n539_));
  INV_X1    g338(.A(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT36), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT78), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT78), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n538_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT79), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT80), .A4(KEYINPUT37), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n534_), .A2(new_n537_), .B1(KEYINPUT78), .B2(new_n544_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(KEYINPUT79), .A3(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n534_), .A2(new_n537_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n543_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n547_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT80), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564_));
  OR2_X1    g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G57gat), .B(G64gat), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n564_), .B(new_n565_), .C1(new_n568_), .C2(KEYINPUT11), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n568_), .A2(KEYINPUT11), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n479_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n572_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT16), .B(G183gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G211gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n575_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(KEYINPUT17), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n563_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n570_), .B(new_n571_), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n528_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n572_), .A2(new_n525_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n587_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(KEYINPUT12), .A3(new_n590_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n572_), .A2(new_n525_), .A3(KEYINPUT12), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n594_), .B2(new_n587_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n292_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n211_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT72), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(KEYINPUT72), .A3(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT71), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n599_), .B1(new_n595_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n604_), .B2(new_n595_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n606_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT73), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n502_), .A2(new_n586_), .A3(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n444_), .B(KEYINPUT109), .Z(new_n614_));
  NOR3_X1   g413(.A1(new_n613_), .A2(G1gat), .A3(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n433_), .A2(new_n441_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n617_), .A2(new_n453_), .A3(new_n446_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n411_), .B1(new_n376_), .B2(new_n410_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n416_), .A2(KEYINPUT104), .A3(new_n421_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n449_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n247_), .A2(new_n421_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n444_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT108), .B1(new_n617_), .B2(new_n453_), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n457_), .B(new_n424_), .C1(new_n433_), .C2(new_n441_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n545_), .A2(new_n550_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n585_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n628_), .A2(new_n630_), .A3(new_n611_), .A4(new_n500_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n451_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n615_), .A2(KEYINPUT38), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n616_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  AND3_X1   g433(.A1(new_n502_), .A2(new_n586_), .A3(new_n612_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT110), .ZN(new_n636_));
  INV_X1    g435(.A(new_n473_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n458_), .A2(new_n459_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .A4(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n502_), .A2(new_n612_), .A3(new_n639_), .A4(new_n586_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT110), .B1(new_n641_), .B2(new_n473_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G8gat), .B1(new_n631_), .B2(new_n638_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT111), .B(KEYINPUT39), .Z(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(KEYINPUT40), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  OAI21_X1  g450(.A(G15gat), .B1(new_n631_), .B2(new_n449_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT41), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n613_), .A2(G15gat), .A3(new_n449_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1326gat));
  OR3_X1    g454(.A1(new_n613_), .A2(G22gat), .A3(new_n421_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G22gat), .B1(new_n631_), .B2(new_n421_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT112), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT112), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n659_), .B(G22gat), .C1(new_n631_), .C2(new_n421_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(KEYINPUT42), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT42), .B1(new_n658_), .B2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT113), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT113), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(new_n656_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n563_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT114), .B1(new_n558_), .B2(new_n562_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n549_), .A2(new_n551_), .B1(new_n556_), .B2(new_n553_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT37), .B1(new_n629_), .B2(KEYINPUT80), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT114), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n448_), .B2(new_n460_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n670_), .B1(new_n677_), .B2(KEYINPUT43), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n584_), .B(new_n501_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT115), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT115), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n671_), .A2(new_n675_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n668_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n683_), .B(new_n679_), .C1(new_n686_), .C2(new_n670_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n681_), .A2(new_n682_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(new_n670_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n680_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n614_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(G29gat), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(G29gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n628_), .A2(new_n629_), .A3(new_n679_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT116), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT116), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n628_), .A2(new_n697_), .A3(new_n679_), .A4(new_n629_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n699_), .B2(new_n451_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n693_), .A2(KEYINPUT117), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT117), .B1(new_n693_), .B2(new_n700_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1328gat));
  AOI21_X1  g502(.A(new_n638_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n688_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  INV_X1    g505(.A(G36gat), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n696_), .A2(new_n707_), .A3(new_n639_), .A4(new_n698_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(KEYINPUT46), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n707_), .B1(new_n688_), .B2(new_n704_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n708_), .B(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n710_), .A2(new_n715_), .ZN(G1329gat));
  AOI21_X1  g515(.A(new_n449_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n688_), .A2(G43gat), .A3(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(KEYINPUT118), .B(G43gat), .Z(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n699_), .B2(new_n449_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT47), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n723_), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1330gat));
  AOI21_X1  g524(.A(new_n421_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n688_), .A2(G50gat), .A3(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n464_), .B1(new_n699_), .B2(new_n421_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1331gat));
  NOR2_X1   g528(.A1(new_n461_), .A2(new_n500_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n611_), .B(KEYINPUT73), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n630_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n451_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n611_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n735_), .A3(new_n586_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(new_n614_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n734_), .B1(new_n737_), .B2(new_n733_), .ZN(G1332gat));
  OAI21_X1  g537(.A(G64gat), .B1(new_n732_), .B2(new_n638_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT48), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n638_), .A2(G64gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT119), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n736_), .B2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n732_), .B2(new_n449_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT49), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n736_), .A2(G71gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n449_), .B2(new_n746_), .ZN(G1334gat));
  OR3_X1    g546(.A1(new_n736_), .A2(G78gat), .A3(new_n421_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G78gat), .B1(new_n732_), .B2(new_n421_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT120), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(G78gat), .C1(new_n732_), .C2(new_n421_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n750_), .A2(KEYINPUT50), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT50), .B1(new_n750_), .B2(new_n752_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n748_), .B1(new_n753_), .B2(new_n754_), .ZN(G1335gat));
  INV_X1    g554(.A(G85gat), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n731_), .A2(new_n629_), .A3(new_n628_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n500_), .A2(new_n584_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n759_), .B2(new_n614_), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n685_), .A2(new_n668_), .B1(new_n461_), .B2(new_n669_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n735_), .A3(new_n758_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(new_n756_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n763_), .B2(new_n451_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT121), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT121), .B(new_n760_), .C1(new_n763_), .C2(new_n451_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1336gat));
  INV_X1    g567(.A(G92gat), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n762_), .A2(new_n769_), .A3(new_n638_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n759_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n639_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n769_), .B2(new_n772_), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n513_), .A3(new_n247_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G99gat), .B1(new_n762_), .B2(new_n449_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n771_), .A2(new_n514_), .A3(new_n410_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n761_), .A2(new_n735_), .A3(new_n410_), .A4(new_n758_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT55), .B1(new_n594_), .B2(new_n587_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n587_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n594_), .B2(KEYINPUT55), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n794_), .B(new_n791_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n789_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n788_), .B1(new_n796_), .B2(new_n599_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n599_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n793_), .A2(new_n795_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT56), .B(new_n798_), .C1(new_n799_), .C2(new_n789_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n482_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n487_), .A2(new_n483_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n495_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n497_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(new_n603_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n603_), .A4(new_n806_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n563_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n602_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n500_), .B1(new_n812_), .B2(new_n600_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n805_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n560_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT57), .B(new_n560_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n811_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n611_), .A2(new_n586_), .A3(new_n501_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT54), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n611_), .A2(new_n586_), .A3(new_n823_), .A4(new_n501_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n820_), .A2(new_n585_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n639_), .A2(new_n614_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n623_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n500_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n820_), .A2(new_n585_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n822_), .A2(new_n824_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n450_), .A4(new_n826_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n623_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n836_), .A2(new_n833_), .A3(new_n837_), .A4(new_n826_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n835_), .A2(new_n500_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n829_), .B1(new_n839_), .B2(G113gat), .ZN(G1340gat));
  NAND3_X1  g639(.A1(new_n835_), .A2(new_n731_), .A3(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G120gat), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(KEYINPUT60), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n611_), .B2(KEYINPUT60), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n836_), .A2(new_n826_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(new_n848_), .ZN(G1341gat));
  AOI21_X1  g648(.A(G127gat), .B1(new_n828_), .B2(new_n584_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n835_), .A2(new_n838_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n584_), .A2(G127gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1342gat));
  NAND4_X1  g652(.A1(new_n835_), .A2(G134gat), .A3(new_n563_), .A4(new_n838_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n828_), .A2(new_n629_), .ZN(new_n855_));
  INV_X1    g654(.A(G134gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n854_), .A2(new_n857_), .ZN(G1343gat));
  NOR4_X1   g657(.A1(new_n825_), .A2(new_n247_), .A3(new_n421_), .A4(new_n827_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n500_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n731_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n584_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n859_), .B2(new_n629_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n684_), .A2(new_n540_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n859_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n639_), .A2(new_n614_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n825_), .A2(new_n623_), .A3(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(KEYINPUT125), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n825_), .A2(new_n873_), .A3(new_n623_), .A4(new_n870_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n330_), .B(new_n500_), .C1(new_n872_), .C2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n871_), .A2(new_n500_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(G169gat), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT62), .B(new_n210_), .C1(new_n871_), .C2(new_n500_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(G1348gat));
  INV_X1    g679(.A(new_n870_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n836_), .A2(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n882_), .A2(new_n211_), .A3(new_n612_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n735_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n223_), .ZN(G1349gat));
  AOI21_X1  g684(.A(G183gat), .B1(new_n871_), .B2(new_n584_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n874_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n873_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n585_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n214_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n889_), .B2(new_n890_), .ZN(G1350gat));
  OAI211_X1 g690(.A(new_n629_), .B(new_n215_), .C1(new_n872_), .C2(new_n874_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n887_), .A2(new_n888_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n893_));
  INV_X1    g692(.A(G190gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1351gat));
  INV_X1    g694(.A(new_n446_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n825_), .A2(new_n638_), .A3(new_n247_), .A4(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n500_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g698(.A(new_n247_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n900_), .A2(new_n639_), .A3(new_n446_), .A4(new_n731_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n297_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT127), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n897_), .A2(new_n904_), .A3(new_n297_), .A4(new_n731_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n897_), .A2(new_n907_), .A3(new_n731_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(G204gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n910_), .ZN(G1353gat));
  NAND2_X1  g710(.A1(new_n897_), .A2(new_n584_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT63), .B(G211gat), .Z(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n912_), .B2(new_n914_), .ZN(G1354gat));
  AOI21_X1  g714(.A(G218gat), .B1(new_n897_), .B2(new_n629_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n897_), .A2(new_n563_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(G218gat), .B2(new_n917_), .ZN(G1355gat));
endmodule


