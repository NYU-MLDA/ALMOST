//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n213_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n212_), .A2(new_n218_), .A3(KEYINPUT86), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224_));
  XOR2_X1   g023(.A(G113gat), .B(G120gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT1), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n216_), .A2(new_n230_), .A3(new_n217_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n213_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT85), .ZN(new_n234_));
  XOR2_X1   g033(.A(G141gat), .B(G148gat), .Z(new_n235_));
  AND3_X1   g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n223_), .B(new_n226_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT97), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n235_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT85), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n226_), .B1(new_n243_), .B2(new_n223_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n223_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT97), .ZN(new_n247_));
  INV_X1    g046(.A(new_n226_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n202_), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n248_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT97), .A3(new_n238_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(new_n249_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n202_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n253_), .B2(KEYINPUT4), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n251_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G1gat), .B(G29gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT98), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G57gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n251_), .B(new_n263_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT94), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n271_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT25), .B(G183gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT26), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G190gat), .ZN(new_n279_));
  INV_X1    g078(.A(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT26), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT24), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT93), .B1(new_n284_), .B2(KEYINPUT24), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n269_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n268_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n288_), .A2(new_n269_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n286_), .B2(new_n285_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(KEYINPUT94), .A3(new_n276_), .A4(new_n282_), .ZN(new_n293_));
  INV_X1    g092(.A(G183gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n280_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n274_), .A2(new_n275_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT22), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G169gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT22), .ZN(new_n300_));
  INV_X1    g099(.A(G176gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n284_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT95), .A2(G169gat), .A3(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n302_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT96), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n296_), .A2(new_n302_), .A3(new_n306_), .A4(KEYINPUT96), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n290_), .A2(new_n293_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(G197gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(G204gat), .ZN(new_n314_));
  INV_X1    g113(.A(G204gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(G197gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT21), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G211gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(G218gat), .ZN(new_n319_));
  INV_X1    g118(.A(G218gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(G211gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT88), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n313_), .B2(G204gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n313_), .A2(G204gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n315_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n317_), .B(new_n322_), .C1(new_n327_), .C2(KEYINPUT21), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT89), .B1(new_n319_), .B2(new_n321_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(G211gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n318_), .A2(G218gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT89), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n327_), .A3(KEYINPUT21), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n312_), .A2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n328_), .A2(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT22), .B1(new_n299_), .B2(KEYINPUT79), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n301_), .C1(KEYINPUT79), .C2(new_n298_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(new_n284_), .A3(new_n296_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT26), .B1(new_n341_), .B2(new_n280_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n278_), .A2(KEYINPUT75), .A3(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n277_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n277_), .A2(KEYINPUT76), .A3(new_n342_), .A4(new_n343_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n271_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT77), .B1(new_n285_), .B2(new_n269_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n299_), .A2(new_n301_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT24), .A4(new_n284_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n271_), .A2(new_n274_), .A3(KEYINPUT78), .A4(new_n275_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n351_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n337_), .B(new_n340_), .C1(new_n348_), .C2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n336_), .A2(KEYINPUT20), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n340_), .B1(new_n348_), .B2(new_n358_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(new_n335_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n362_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n337_), .A2(new_n290_), .A3(new_n293_), .A4(new_n311_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT18), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  AND2_X1   g172(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT99), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT99), .ZN(new_n376_));
  INV_X1    g175(.A(new_n373_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AND4_X1   g178(.A1(new_n363_), .A2(new_n369_), .A3(new_n375_), .A4(new_n379_), .ZN(new_n380_));
  AND4_X1   g179(.A1(KEYINPUT20), .A2(new_n336_), .A3(new_n367_), .A4(new_n359_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n337_), .A2(KEYINPUT91), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n292_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT91), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n335_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n382_), .A2(new_n307_), .A3(new_n383_), .A4(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n367_), .B1(new_n366_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n374_), .B1(new_n381_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT100), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT100), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n390_), .B(new_n374_), .C1(new_n381_), .C2(new_n387_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n380_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n267_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n266_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n264_), .A2(new_n394_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n251_), .B(new_n396_), .C1(new_n255_), .C2(new_n257_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n363_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n373_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n254_), .A2(new_n249_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n263_), .B1(new_n401_), .B2(new_n256_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n202_), .B1(new_n253_), .B2(KEYINPUT4), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n255_), .B2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n395_), .A2(new_n397_), .A3(new_n400_), .A4(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G228gat), .ZN(new_n406_));
  INV_X1    g205(.A(G233gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT29), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n243_), .B2(new_n223_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n335_), .B(KEYINPUT91), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n408_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n246_), .A2(KEYINPUT29), .ZN(new_n413_));
  INV_X1    g212(.A(new_n408_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n335_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT90), .B1(new_n413_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n418_));
  AOI211_X1 g217(.A(new_n418_), .B(new_n415_), .C1(new_n246_), .C2(KEYINPUT29), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n412_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(new_n412_), .C1(new_n417_), .C2(new_n419_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n243_), .A2(new_n409_), .A3(new_n223_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n426_));
  XOR2_X1   g225(.A(G22gat), .B(G50gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n425_), .B(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n422_), .A2(KEYINPUT92), .A3(new_n424_), .A4(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT92), .B1(new_n420_), .B2(new_n421_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n418_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n413_), .A2(KEYINPUT90), .A3(new_n416_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n423_), .B1(new_n435_), .B2(new_n412_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n424_), .ZN(new_n437_));
  OAI22_X1  g236(.A1(new_n431_), .A2(new_n432_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n393_), .A2(new_n405_), .A3(new_n430_), .A4(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(KEYINPUT81), .B(G15gat), .Z(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  INV_X1    g245(.A(new_n340_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n351_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n346_), .A2(new_n347_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G43gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n450_), .A2(new_n452_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n454_), .A2(new_n248_), .A3(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n450_), .A2(new_n452_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n226_), .B1(new_n457_), .B2(new_n453_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n446_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n248_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n453_), .A3(new_n226_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n444_), .B(new_n445_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n459_), .A2(KEYINPUT83), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT83), .B1(new_n459_), .B2(new_n463_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n438_), .A2(new_n430_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT27), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n468_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n377_), .B1(new_n381_), .B2(new_n387_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n363_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT27), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n265_), .A3(new_n266_), .A4(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n466_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n472_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n467_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n459_), .A2(new_n463_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n267_), .A2(new_n477_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n439_), .A2(new_n474_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT70), .ZN(new_n483_));
  INV_X1    g282(.A(G36gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(G29gat), .ZN(new_n485_));
  INV_X1    g284(.A(G29gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G36gat), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n485_), .A2(new_n487_), .A3(KEYINPUT70), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n487_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n482_), .A2(KEYINPUT70), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n480_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G1gat), .A2(G8gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT14), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G8gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n495_), .A2(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n495_), .B(new_n503_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n506_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n504_), .A2(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G113gat), .B(G141gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(G169gat), .B(G197gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n514_), .A2(KEYINPUT74), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(KEYINPUT74), .ZN(new_n516_));
  OAI22_X1  g315(.A1(new_n515_), .A2(new_n516_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G85gat), .B(G92gat), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT10), .B(G99gat), .Z(new_n520_));
  INV_X1    g319(.A(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT6), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(G99gat), .A3(G106gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT64), .B(G92gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT9), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(G85gat), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n519_), .A2(new_n522_), .A3(new_n527_), .A4(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n533_), .B(new_n534_), .C1(G99gat), .C2(G106gat), .ZN(new_n535_));
  INV_X1    g334(.A(G99gat), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(new_n521_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n527_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT66), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT66), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n541_), .A3(new_n527_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT8), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n518_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n527_), .A2(KEYINPUT67), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n524_), .A2(new_n526_), .A3(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n550_), .A3(new_n538_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n518_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT8), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n532_), .B1(new_n547_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n557_));
  XOR2_X1   g356(.A(G71gat), .B(G78gat), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OR3_X1    g360(.A1(new_n554_), .A2(KEYINPUT12), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n545_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n544_), .B1(new_n551_), .B2(new_n518_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n531_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n531_), .B(new_n561_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT12), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n567_), .A2(new_n568_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n571_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n562_), .A2(new_n569_), .B1(G230gat), .B2(G233gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n582_), .B2(new_n574_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n581_), .A2(new_n583_), .A3(KEYINPUT13), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT13), .B1(new_n581_), .B2(new_n583_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT68), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n580_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n582_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(new_n583_), .A3(KEYINPUT13), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT68), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n517_), .B1(new_n587_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n479_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n489_), .A2(new_n494_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n531_), .B(new_n596_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT34), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(KEYINPUT71), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n601_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n495_), .B(KEYINPUT15), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n554_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n597_), .A2(new_n603_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n604_), .B(new_n606_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n597_), .A2(new_n603_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n497_), .A2(new_n565_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n611_), .B(new_n612_), .C1(KEYINPUT71), .C2(new_n605_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n610_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n616_), .B(KEYINPUT36), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT72), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT37), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  NOR4_X1   g424(.A1(new_n618_), .A2(new_n621_), .A3(KEYINPUT72), .A4(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n561_), .B(new_n503_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G127gat), .B(G155gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n630_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n638_), .B1(new_n636_), .B2(new_n630_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT73), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n627_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n267_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(G1gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n595_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(KEYINPUT38), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n594_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT102), .B(new_n517_), .C1(new_n587_), .C2(new_n593_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n622_), .B(KEYINPUT103), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n479_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n653_), .A2(new_n640_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n643_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT38), .B1(new_n647_), .B2(new_n648_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT104), .B(KEYINPUT38), .C1(new_n647_), .C2(new_n648_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n658_), .B(KEYINPUT105), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1324gat));
  XNOR2_X1  g466(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n653_), .A2(new_n640_), .A3(new_n475_), .A4(new_n655_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G8gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n595_), .A2(new_n642_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G8gat), .B1(new_n469_), .B2(new_n472_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n674_), .A2(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n673_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n668_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n673_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT106), .B1(new_n669_), .B2(G8gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n675_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n677_), .A2(new_n678_), .ZN(new_n686_));
  AND4_X1   g485(.A1(new_n681_), .A2(new_n685_), .A3(new_n686_), .A4(new_n668_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n682_), .A2(new_n687_), .ZN(G1325gat));
  INV_X1    g487(.A(new_n466_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n676_), .A2(G15gat), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n656_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n466_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT41), .B1(new_n692_), .B2(G15gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n467_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(G22gat), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G22gat), .ZN(new_n699_));
  INV_X1    g498(.A(new_n467_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(G22gat), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT110), .Z(new_n702_));
  OAI22_X1  g501(.A1(new_n698_), .A2(new_n699_), .B1(new_n676_), .B2(new_n702_), .ZN(G1327gat));
  INV_X1    g502(.A(new_n622_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n640_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n595_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G29gat), .B1(new_n707_), .B2(new_n267_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT111), .B1(new_n624_), .B2(new_n626_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n621_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n610_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n623_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n625_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n622_), .A2(new_n623_), .A3(KEYINPUT37), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n710_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n479_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n479_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n439_), .A2(new_n474_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n476_), .A2(new_n478_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n627_), .A2(KEYINPUT43), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n721_), .A2(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n640_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n653_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n709_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(new_n726_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n710_), .A2(new_n717_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n725_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT112), .B1(new_n733_), .B2(KEYINPUT43), .ZN(new_n734_));
  INV_X1    g533(.A(new_n722_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n729_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(KEYINPUT44), .A3(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n730_), .A2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n643_), .A2(new_n486_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n708_), .B1(new_n739_), .B2(new_n740_), .ZN(G1328gat));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n730_), .A2(new_n738_), .A3(new_n475_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G36gat), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n595_), .A2(new_n484_), .A3(new_n475_), .A4(new_n705_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT45), .Z(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n744_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n742_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n746_), .B(new_n749_), .C1(new_n743_), .C2(G36gat), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1329gat));
  INV_X1    g550(.A(new_n477_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n730_), .A2(new_n738_), .A3(G43gat), .A4(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(G43gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n706_), .B2(new_n689_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT47), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1330gat));
  AOI21_X1  g560(.A(G50gat), .B1(new_n707_), .B2(new_n467_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n467_), .A2(G50gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n739_), .B2(new_n763_), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n584_), .A2(new_n585_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT68), .ZN(new_n766_));
  INV_X1    g565(.A(new_n593_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n517_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n640_), .ZN(new_n770_));
  NOR4_X1   g569(.A1(new_n768_), .A2(new_n479_), .A3(new_n654_), .A4(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G57gat), .B1(new_n772_), .B2(new_n643_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n768_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT115), .A3(new_n642_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n479_), .A2(new_n517_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n768_), .B2(new_n641_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT116), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n643_), .A2(G57gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n773_), .B1(new_n780_), .B2(new_n781_), .ZN(G1332gat));
  INV_X1    g581(.A(G64gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n771_), .B2(new_n475_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT48), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n475_), .A2(new_n783_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n780_), .B2(new_n786_), .ZN(G1333gat));
  NOR3_X1   g586(.A1(new_n780_), .A2(G71gat), .A3(new_n689_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n771_), .A2(new_n466_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G71gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G71gat), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n788_), .A2(KEYINPUT117), .A3(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT117), .B1(new_n788_), .B2(new_n793_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1334gat));
  INV_X1    g595(.A(G78gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n771_), .B2(new_n467_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT50), .Z(new_n799_));
  NAND2_X1  g598(.A1(new_n467_), .A2(new_n797_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n780_), .B2(new_n800_), .ZN(G1335gat));
  INV_X1    g600(.A(G85gat), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n768_), .A2(new_n640_), .A3(new_n517_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n721_), .A2(new_n722_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n731_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n802_), .B1(new_n808_), .B2(new_n267_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n776_), .A2(new_n774_), .A3(new_n705_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n643_), .A2(G85gat), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n809_), .A2(new_n812_), .ZN(G1336gat));
  INV_X1    g612(.A(new_n810_), .ZN(new_n814_));
  AOI21_X1  g613(.A(G92gat), .B1(new_n814_), .B2(new_n475_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT119), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n475_), .A2(new_n528_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n808_), .B2(new_n817_), .ZN(G1337gat));
  AOI21_X1  g617(.A(new_n536_), .B1(new_n806_), .B2(new_n466_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n814_), .A2(new_n520_), .A3(new_n752_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n819_), .A2(new_n820_), .B1(KEYINPUT120), .B2(KEYINPUT51), .ZN(new_n821_));
  NAND2_X1  g620(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1338gat));
  NAND3_X1  g622(.A1(new_n814_), .A2(new_n521_), .A3(new_n467_), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT52), .B(new_n521_), .C1(new_n806_), .C2(new_n467_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n736_), .A2(new_n467_), .A3(new_n803_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(G106gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT53), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n824_), .C1(new_n825_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1339gat));
  NAND3_X1  g632(.A1(new_n476_), .A2(new_n267_), .A3(new_n752_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT122), .Z(new_n835_));
  OR2_X1    g634(.A1(new_n514_), .A2(KEYINPUT74), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n514_), .A2(KEYINPUT74), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n504_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n513_), .B1(new_n508_), .B2(new_n506_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n836_), .A2(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n581_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n582_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n571_), .B2(new_n570_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n580_), .B1(new_n582_), .B2(new_n842_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n844_), .A2(KEYINPUT56), .A3(new_n845_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n850_), .A2(KEYINPUT58), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n627_), .B1(new_n850_), .B2(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n517_), .A2(new_n581_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n581_), .A2(new_n583_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n840_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n704_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n851_), .A2(new_n852_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n857_), .A2(new_n858_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n640_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n627_), .A2(new_n640_), .A3(new_n769_), .A4(new_n765_), .ZN(new_n862_));
  OR2_X1    g661(.A1(KEYINPUT121), .A2(KEYINPUT54), .ZN(new_n863_));
  NAND2_X1  g662(.A1(KEYINPUT121), .A2(KEYINPUT54), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n835_), .B1(new_n861_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G113gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n517_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n861_), .A2(new_n866_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n867_), .B(new_n871_), .C1(new_n872_), .C2(KEYINPUT123), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  OAI221_X1 g673(.A(new_n835_), .B1(new_n874_), .B2(KEYINPUT59), .C1(new_n861_), .C2(new_n866_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n769_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n870_), .B1(new_n876_), .B2(new_n869_), .ZN(G1340gat));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n768_), .B2(KEYINPUT60), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n868_), .B(new_n879_), .C1(KEYINPUT60), .C2(new_n878_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n768_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n878_), .ZN(G1341gat));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n868_), .A2(new_n883_), .A3(new_n640_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n728_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(G1342gat));
  AOI21_X1  g685(.A(G134gat), .B1(new_n868_), .B2(new_n654_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n873_), .A2(new_n875_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT124), .B(G134gat), .Z(new_n889_));
  NOR2_X1   g688(.A1(new_n627_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n888_), .B2(new_n890_), .ZN(G1343gat));
  OR2_X1    g690(.A1(new_n861_), .A2(new_n866_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n700_), .A2(new_n466_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n894_), .A2(new_n643_), .A3(new_n475_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n517_), .A3(new_n895_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT125), .B(G141gat), .Z(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n892_), .A2(new_n774_), .A3(new_n895_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n892_), .A2(new_n640_), .A3(new_n895_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  AND2_X1   g702(.A1(new_n892_), .A2(new_n895_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n654_), .ZN(new_n905_));
  INV_X1    g704(.A(G162gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n718_), .A2(new_n906_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n905_), .A2(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n643_), .A2(new_n475_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n689_), .A2(new_n467_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n872_), .A2(new_n769_), .A3(new_n910_), .A4(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n909_), .B1(new_n913_), .B2(new_n299_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n910_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n892_), .A2(new_n517_), .A3(new_n916_), .A4(new_n911_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n914_), .A2(new_n915_), .A3(new_n918_), .ZN(G1348gat));
  NAND4_X1  g718(.A1(new_n892_), .A2(new_n774_), .A3(new_n916_), .A4(new_n911_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT126), .B(G176gat), .Z(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n872_), .A2(new_n910_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n301_), .A2(KEYINPUT126), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n923_), .A2(new_n774_), .A3(new_n911_), .A4(new_n924_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n922_), .A2(new_n925_), .ZN(G1349gat));
  NAND4_X1  g725(.A1(new_n892_), .A2(new_n640_), .A3(new_n916_), .A4(new_n911_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n927_), .A2(new_n294_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n277_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1350gat));
  NAND2_X1  g729(.A1(new_n892_), .A2(new_n916_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n931_), .A2(new_n627_), .A3(new_n912_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n923_), .A2(new_n911_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n654_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n932_), .A2(new_n280_), .B1(new_n933_), .B2(new_n934_), .ZN(G1351gat));
  NAND4_X1  g734(.A1(new_n892_), .A2(new_n517_), .A3(new_n893_), .A4(new_n916_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  XNOR2_X1  g736(.A(KEYINPUT127), .B(G204gat), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n923_), .A2(new_n774_), .A3(new_n893_), .A4(new_n938_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n931_), .A2(new_n768_), .A3(new_n894_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1353gat));
  AOI21_X1  g741(.A(new_n728_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n892_), .A2(new_n893_), .A3(new_n916_), .A4(new_n943_), .ZN(new_n944_));
  OR2_X1    g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1354gat));
  NAND4_X1  g745(.A1(new_n923_), .A2(new_n320_), .A3(new_n654_), .A4(new_n893_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n931_), .A2(new_n627_), .A3(new_n894_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n948_), .B2(new_n320_), .ZN(G1355gat));
endmodule


