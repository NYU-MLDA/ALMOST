//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G204gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G197gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(new_n207_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT21), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G211gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(G218gat), .ZN(new_n217_));
  INV_X1    g016(.A(G218gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(G211gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT89), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(G211gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(G218gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT89), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n213_), .A2(new_n210_), .A3(KEYINPUT88), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n213_), .A2(new_n210_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(KEYINPUT21), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n215_), .A2(new_n225_), .A3(new_n227_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT90), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n223_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n220_), .A2(KEYINPUT90), .A3(new_n224_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(KEYINPUT21), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT91), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n236_), .A2(new_n237_), .A3(new_n242_), .A4(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n232_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT25), .B(G183gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT94), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT26), .B(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT95), .A3(KEYINPUT24), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(KEYINPUT24), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT95), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n247_), .A2(new_n248_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(KEYINPUT23), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT82), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n256_), .B(KEYINPUT23), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(KEYINPUT82), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT24), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n251_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(G183gat), .B2(G190gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n249_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT22), .B(G169gat), .ZN(new_n265_));
  INV_X1    g064(.A(G176gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n255_), .A2(new_n262_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT20), .B1(new_n244_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n238_), .B1(new_n225_), .B2(new_n233_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n242_), .B1(new_n270_), .B2(new_n237_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n243_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n231_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT22), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G169gat), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n277_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT81), .B1(new_n277_), .B2(KEYINPUT22), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n276_), .A2(new_n278_), .A3(new_n266_), .A4(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n280_), .A2(new_n249_), .ZN(new_n281_));
  OAI221_X1 g080(.A(new_n258_), .B1(G183gat), .B2(G190gat), .C1(new_n259_), .C2(KEYINPUT82), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n252_), .A2(new_n251_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n251_), .A2(new_n261_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n283_), .A2(new_n259_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT26), .ZN(new_n286_));
  OR3_X1    g085(.A1(new_n286_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(G190gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT79), .B1(new_n286_), .B2(G190gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n287_), .A2(new_n245_), .A3(new_n288_), .A4(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n281_), .A2(new_n282_), .B1(new_n285_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n273_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n269_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n244_), .B2(new_n268_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT96), .B1(new_n273_), .B2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT96), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n244_), .A2(new_n300_), .A3(new_n291_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n295_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n296_), .B1(new_n303_), .B2(KEYINPUT99), .ZN(new_n304_));
  INV_X1    g103(.A(new_n295_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n273_), .A2(KEYINPUT96), .A3(new_n292_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n300_), .B1(new_n244_), .B2(new_n291_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI211_X1 g107(.A(KEYINPUT99), .B(new_n305_), .C1(new_n308_), .C2(new_n298_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n206_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n311_));
  AOI211_X1 g110(.A(new_n297_), .B(new_n295_), .C1(new_n244_), .C2(new_n268_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT97), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n295_), .B1(new_n269_), .B2(new_n293_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n308_), .A2(KEYINPUT97), .A3(new_n312_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n315_), .A2(new_n206_), .A3(new_n316_), .A4(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT27), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n202_), .B1(new_n311_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n206_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n305_), .B1(new_n308_), .B2(new_n298_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT99), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n269_), .A2(new_n293_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n322_), .A2(new_n323_), .B1(new_n295_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n321_), .B1(new_n325_), .B2(new_n309_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n326_), .A2(KEYINPUT101), .A3(KEYINPUT27), .A4(new_n318_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n320_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n329_));
  NOR2_X1   g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT84), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT3), .Z(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT2), .Z(new_n336_));
  OAI211_X1 g135(.A(new_n331_), .B(new_n332_), .C1(new_n334_), .C2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n332_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n331_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n333_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n335_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n329_), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  INV_X1    g144(.A(new_n329_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n337_), .A2(new_n342_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G22gat), .B(G50gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G233gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n351_), .A2(KEYINPUT86), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(KEYINPUT86), .ZN(new_n353_));
  OAI21_X1  g152(.A(G228gat), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n343_), .A2(KEYINPUT29), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n355_), .B1(new_n357_), .B2(new_n244_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n273_), .A2(new_n356_), .A3(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n350_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n350_), .B(new_n364_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT93), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n350_), .A2(new_n364_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(KEYINPUT92), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .A4(new_n369_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n365_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n317_), .A2(new_n316_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT97), .B1(new_n308_), .B2(new_n312_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n321_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT27), .B1(new_n379_), .B2(new_n318_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(G127gat), .B(G134gat), .Z(new_n383_));
  XOR2_X1   g182(.A(G113gat), .B(G120gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n343_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n337_), .A2(new_n342_), .A3(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT4), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n343_), .A2(new_n390_), .A3(new_n386_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n382_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G85gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT0), .B(G57gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n387_), .A2(new_n388_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n382_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n393_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n397_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n399_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(new_n392_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G15gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT30), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n291_), .B(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT83), .B1(new_n386_), .B2(KEYINPUT31), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(KEYINPUT31), .B2(new_n386_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n410_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n413_), .B(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n406_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n328_), .A2(new_n376_), .A3(new_n381_), .A4(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n376_), .A2(new_n380_), .A3(new_n406_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n315_), .A2(new_n420_), .A3(new_n316_), .A4(new_n317_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n404_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n379_), .A2(new_n318_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n403_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n397_), .B1(new_n398_), .B2(new_n382_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT98), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(KEYINPUT98), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n389_), .A2(new_n382_), .A3(new_n391_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n403_), .A2(new_n425_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n426_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n421_), .A2(new_n423_), .B1(new_n424_), .B2(new_n433_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n419_), .A2(new_n328_), .B1(new_n376_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n416_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n418_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT72), .B(G8gat), .ZN(new_n438_));
  INV_X1    g237(.A(G1gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G15gat), .B(G22gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G1gat), .B(G8gat), .Z(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G29gat), .B(G36gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT69), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G43gat), .B(G50gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G229gat), .A2(G233gat), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n446_), .A2(new_n447_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n452_), .B(KEYINPUT15), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n455_), .A2(KEYINPUT76), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT76), .B1(new_n455_), .B2(new_n456_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n453_), .B(new_n454_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n448_), .B(new_n452_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n454_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G169gat), .B(G197gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT77), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n459_), .A2(new_n468_), .A3(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT78), .B1(new_n470_), .B2(new_n471_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n437_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n479_));
  INV_X1    g278(.A(G231gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(new_n351_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n448_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT67), .B(G71gat), .ZN(new_n483_));
  INV_X1    g282(.A(G78gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n488_), .B1(new_n491_), .B2(new_n485_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n446_), .B(new_n447_), .C1(new_n480_), .C2(new_n351_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n482_), .B2(new_n494_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G127gat), .B(G155gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n482_), .A2(new_n494_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n492_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(new_n499_), .A3(new_n495_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n502_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G183gat), .B(G211gat), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n504_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n479_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n504_), .A2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n498_), .A2(new_n479_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT34), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT10), .B(G99gat), .Z(new_n523_));
  INV_X1    g322(.A(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT65), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G85gat), .B(G92gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT9), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(G85gat), .A3(G92gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT6), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n526_), .A2(new_n529_), .A3(new_n531_), .A4(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT7), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n535_), .B1(new_n540_), .B2(new_n528_), .ZN(new_n541_));
  AOI211_X1 g340(.A(KEYINPUT8), .B(new_n527_), .C1(new_n538_), .C2(new_n533_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n534_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n456_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n522_), .B1(new_n544_), .B2(KEYINPUT70), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n452_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G190gat), .B(G218gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT71), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n546_), .A2(new_n549_), .B1(KEYINPUT36), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n549_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n545_), .B2(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n555_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n560_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n558_), .A2(new_n545_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n565_), .B(new_n553_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n555_), .A2(new_n560_), .A3(new_n557_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT64), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n543_), .A2(new_n492_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n493_), .B(new_n534_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(KEYINPUT12), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n543_), .A2(new_n578_), .A3(new_n492_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n574_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n576_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n574_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G120gat), .B(G148gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n582_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n588_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT13), .B1(new_n589_), .B2(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n519_), .A2(new_n571_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n478_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n406_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n596_), .A2(G1gat), .A3(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT38), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT102), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n561_), .A2(new_n562_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n593_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n472_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND4_X1   g404(.A1(new_n437_), .A2(new_n519_), .A3(new_n602_), .A4(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n439_), .B1(new_n606_), .B2(new_n406_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n598_), .B2(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(G8gat), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n328_), .A2(new_n381_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT39), .Z(new_n613_));
  INV_X1    g412(.A(new_n596_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n611_), .A3(new_n438_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n606_), .B2(new_n436_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT41), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(new_n618_), .A3(new_n436_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT103), .ZN(G1326gat));
  INV_X1    g422(.A(G22gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n376_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n606_), .B2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT42), .Z(new_n627_));
  NOR2_X1   g426(.A1(new_n376_), .A2(G22gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT104), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n596_), .B2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n519_), .ZN(new_n631_));
  AND4_X1   g430(.A1(new_n478_), .A2(new_n631_), .A3(new_n601_), .A4(new_n593_), .ZN(new_n632_));
  INV_X1    g431(.A(G29gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n406_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  INV_X1    g434(.A(new_n571_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n419_), .A2(new_n328_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n434_), .A2(new_n376_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n436_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n418_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n635_), .B(new_n636_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT105), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n437_), .A2(new_n643_), .A3(new_n635_), .A4(new_n636_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT43), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n605_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT106), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n631_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n650_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n651_), .B1(new_n647_), .B2(new_n605_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT44), .B1(new_n655_), .B2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(KEYINPUT107), .A3(new_n406_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT107), .B1(new_n657_), .B2(new_n406_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n634_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n632_), .A2(new_n662_), .A3(new_n611_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT45), .ZN(new_n664_));
  INV_X1    g463(.A(new_n611_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n666_), .B2(new_n662_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT46), .B(new_n664_), .C1(new_n666_), .C2(new_n662_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  INV_X1    g470(.A(KEYINPUT47), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n650_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n652_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n436_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G43gat), .ZN(new_n676_));
  INV_X1    g475(.A(G43gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n632_), .A2(new_n677_), .A3(new_n436_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n672_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n416_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n672_), .B(new_n678_), .C1(new_n680_), .C2(new_n677_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1330gat));
  INV_X1    g482(.A(G50gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n632_), .A2(new_n684_), .A3(new_n625_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n657_), .A2(new_n625_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT108), .B1(new_n686_), .B2(G50gat), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n688_), .B(new_n684_), .C1(new_n657_), .C2(new_n625_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n687_), .B2(new_n689_), .ZN(G1331gat));
  NAND2_X1  g489(.A1(new_n437_), .A2(new_n604_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT109), .ZN(new_n692_));
  AND4_X1   g491(.A1(new_n519_), .A2(new_n692_), .A3(new_n571_), .A4(new_n603_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n406_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n631_), .A2(new_n477_), .A3(new_n593_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n695_), .A2(new_n437_), .A3(new_n602_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(G57gat), .A3(new_n406_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT110), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1332gat));
  INV_X1    g498(.A(G64gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(new_n700_), .A3(new_n611_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n696_), .B2(new_n611_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1333gat));
  INV_X1    g504(.A(G71gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n696_), .B2(new_n436_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT49), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n693_), .A2(new_n706_), .A3(new_n436_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT112), .ZN(G1334gat));
  AOI21_X1  g510(.A(new_n484_), .B1(new_n696_), .B2(new_n625_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT50), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n693_), .A2(new_n484_), .A3(new_n625_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1335gat));
  AND4_X1   g514(.A1(new_n631_), .A2(new_n692_), .A3(new_n601_), .A4(new_n603_), .ZN(new_n716_));
  INV_X1    g515(.A(G85gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n406_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n519_), .A2(new_n593_), .A3(new_n472_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n647_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n597_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1336gat));
  INV_X1    g521(.A(G92gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n716_), .A2(new_n723_), .A3(new_n611_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G92gat), .B1(new_n720_), .B2(new_n665_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1337gat));
  NOR2_X1   g525(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n716_), .A2(new_n436_), .A3(new_n523_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G99gat), .B1(new_n720_), .B2(new_n416_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT114), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n730_), .B(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n716_), .A2(new_n524_), .A3(new_n625_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n647_), .A2(KEYINPUT115), .A3(new_n625_), .A4(new_n719_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(G106gat), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n720_), .B2(new_n376_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n736_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n736_), .B2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n734_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n734_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  NAND4_X1  g545(.A1(new_n519_), .A2(new_n476_), .A3(new_n571_), .A4(new_n593_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT57), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n459_), .A2(new_n468_), .A3(new_n462_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n468_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n590_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n577_), .A2(new_n574_), .A3(new_n579_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT55), .ZN(new_n755_));
  INV_X1    g554(.A(new_n580_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n580_), .A2(KEYINPUT55), .A3(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n587_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n753_), .B1(new_n760_), .B2(KEYINPUT116), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n587_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n587_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n589_), .A2(new_n590_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n453_), .B(new_n461_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n460_), .A2(new_n454_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n466_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n467_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n761_), .A2(new_n767_), .B1(new_n768_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n750_), .B1(new_n774_), .B2(new_n601_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n768_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n470_), .A2(new_n471_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(KEYINPUT57), .A3(new_n602_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n590_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n760_), .B2(KEYINPUT117), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n764_), .A2(new_n765_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT118), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n636_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT118), .B(KEYINPUT58), .C1(new_n783_), .C2(new_n785_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n775_), .B(new_n781_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n519_), .B1(new_n790_), .B2(KEYINPUT119), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n788_), .A2(new_n789_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n775_), .A4(new_n781_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n749_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n611_), .A2(new_n625_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n597_), .A2(new_n416_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT120), .ZN(new_n800_));
  INV_X1    g599(.A(G113gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(KEYINPUT120), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n472_), .A4(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT59), .B1(new_n795_), .B2(new_n798_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n798_), .B(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n790_), .A2(new_n631_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT123), .B(new_n808_), .C1(new_n809_), .C2(new_n749_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n749_), .B1(new_n631_), .B2(new_n790_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n806_), .A2(new_n807_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n804_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n804_), .B2(new_n815_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n476_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n803_), .B1(new_n819_), .B2(new_n801_), .ZN(G1340gat));
  NAND3_X1  g619(.A1(new_n804_), .A2(new_n815_), .A3(new_n603_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n800_), .A2(new_n802_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G120gat), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n593_), .A2(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n822_), .B1(new_n823_), .B2(new_n827_), .ZN(G1341gat));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n800_), .A2(new_n829_), .A3(new_n519_), .A4(new_n802_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n817_), .A2(new_n818_), .A3(new_n631_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n829_), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n800_), .A2(new_n833_), .A3(new_n601_), .A4(new_n802_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n817_), .A2(new_n818_), .A3(new_n571_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n833_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n795_), .A2(new_n436_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n611_), .A2(new_n376_), .A3(new_n597_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n472_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n603_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n837_), .A2(new_n838_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n631_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  OR3_X1    g646(.A1(new_n844_), .A2(G162gat), .A3(new_n602_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G162gat), .B1(new_n844_), .B2(new_n571_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1347gat));
  NAND2_X1  g649(.A1(new_n611_), .A2(new_n417_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n812_), .A2(new_n625_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(G169gat), .B1(new_n853_), .B2(new_n604_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n855_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n265_), .A3(new_n472_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(G1348gat));
  AOI21_X1  g658(.A(G176gat), .B1(new_n852_), .B2(new_n603_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n795_), .A2(new_n625_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n851_), .A2(new_n266_), .A3(new_n593_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(G1349gat));
  NOR2_X1   g662(.A1(new_n631_), .A2(new_n851_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G183gat), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n812_), .A2(new_n625_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n631_), .A2(new_n851_), .A3(new_n247_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n853_), .B2(new_n571_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n852_), .A2(new_n248_), .A3(new_n601_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1351gat));
  NAND3_X1  g670(.A1(new_n611_), .A2(new_n625_), .A3(new_n597_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n837_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n604_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n208_), .ZN(G1352gat));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n593_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n212_), .ZN(G1353gat));
  AOI21_X1  g677(.A(new_n631_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n837_), .A2(new_n873_), .A3(new_n879_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT125), .B(KEYINPUT126), .Z(new_n881_));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n880_), .B(new_n883_), .ZN(G1354gat));
  NOR3_X1   g683(.A1(new_n874_), .A2(new_n218_), .A3(new_n571_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n874_), .A2(new_n602_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G218gat), .B1(new_n886_), .B2(KEYINPUT127), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n874_), .B2(new_n602_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n887_), .B2(new_n889_), .ZN(G1355gat));
endmodule


