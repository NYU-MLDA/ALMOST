//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G232gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n211_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT77), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT9), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n220_), .B2(KEYINPUT65), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n222_), .A3(KEYINPUT9), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n221_), .B(new_n223_), .C1(G106gat), .C2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT6), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT66), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n234_));
  INV_X1    g033(.A(new_n232_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n226_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n232_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n235_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT67), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n225_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G99gat), .A2(G106gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT69), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  INV_X1    g048(.A(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT7), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT68), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n248_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n252_), .B1(G99gat), .B2(G106gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .A4(new_n247_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n245_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n238_), .A2(new_n239_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n254_), .A2(new_n256_), .A3(new_n247_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n257_), .B1(new_n251_), .B2(KEYINPUT7), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT70), .A3(new_n258_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n244_), .B1(new_n267_), .B2(new_n219_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n258_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n237_), .A2(new_n240_), .A3(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n270_), .A2(new_n244_), .A3(new_n219_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n243_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G29gat), .B(G36gat), .Z(new_n273_));
  XOR2_X1   g072(.A(G43gat), .B(G50gat), .Z(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  OAI21_X1  g074(.A(new_n215_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n265_), .A2(KEYINPUT70), .A3(new_n258_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n265_), .B2(new_n258_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n261_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT8), .B1(new_n280_), .B2(new_n220_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(new_n244_), .A3(new_n219_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n242_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n275_), .B(KEYINPUT15), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n277_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n272_), .A2(KEYINPUT75), .A3(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n276_), .B1(new_n288_), .B2(KEYINPUT76), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT76), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n290_), .A3(new_n287_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n213_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n212_), .B(KEYINPUT80), .ZN(new_n293_));
  AOI211_X1 g092(.A(new_n293_), .B(new_n276_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n207_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  OAI221_X1 g099(.A(new_n296_), .B1(new_n298_), .B2(new_n207_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT37), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(KEYINPUT37), .A3(new_n301_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT19), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT94), .B(G204gat), .Z(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(G197gat), .ZN(new_n311_));
  INV_X1    g110(.A(G197gat), .ZN(new_n312_));
  INV_X1    g111(.A(G204gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT21), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n310_), .B2(G197gat), .ZN(new_n316_));
  OAI221_X1 g115(.A(new_n309_), .B1(new_n311_), .B2(new_n314_), .C1(KEYINPUT21), .C2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n309_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(KEYINPUT21), .A3(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT23), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n332_), .A2(KEYINPUT24), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT95), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n329_), .A2(KEYINPUT95), .A3(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n332_), .A2(KEYINPUT24), .A3(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT25), .B(G183gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G190gat), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(new_n323_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(G183gat), .B2(G190gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n331_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n338_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n320_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n329_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(G169gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n345_), .A2(new_n342_), .A3(new_n333_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n317_), .A2(new_n319_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT20), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n308_), .B1(new_n350_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n320_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n308_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT20), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT18), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G64gat), .B(G92gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n360_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT3), .Z(new_n381_));
  NAND2_X1  g180(.A1(G141gat), .A2(G148gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n382_), .B(KEYINPUT2), .Z(new_n383_));
  OAI211_X1 g182(.A(new_n377_), .B(new_n379_), .C1(new_n381_), .C2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n378_), .B1(KEYINPUT1), .B2(new_n377_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(KEYINPUT1), .B2(new_n377_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n380_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n391_), .A2(new_n392_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n395_), .A2(KEYINPUT92), .ZN(new_n396_));
  OR3_X1    g195(.A1(new_n393_), .A2(new_n394_), .A3(new_n390_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(new_n395_), .A3(KEYINPUT92), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n395_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n389_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT96), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n401_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n376_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n399_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(KEYINPUT4), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n405_), .B2(KEYINPUT4), .ZN(new_n411_));
  AOI22_X1  g210(.A1(KEYINPUT97), .A2(new_n408_), .B1(new_n411_), .B2(new_n406_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n408_), .A2(KEYINPUT97), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n372_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n401_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n404_), .A2(new_n399_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT4), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n410_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n406_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n405_), .A2(new_n407_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n376_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT33), .B(new_n376_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n420_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n376_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n426_), .B(new_n427_), .C1(new_n411_), .C2(new_n406_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n421_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n308_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT99), .B1(new_n361_), .B2(KEYINPUT20), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n358_), .B2(new_n357_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n361_), .A2(KEYINPUT99), .A3(KEYINPUT20), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n430_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n350_), .A2(new_n359_), .A3(new_n308_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT32), .B(new_n368_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n360_), .A2(new_n363_), .A3(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT98), .Z(new_n439_));
  NAND3_X1  g238(.A1(new_n429_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n425_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(G15gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT30), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT31), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n357_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n398_), .A2(new_n396_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n357_), .A2(new_n449_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n446_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n445_), .A3(new_n454_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n384_), .A2(new_n388_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT28), .B1(new_n462_), .B2(KEYINPUT29), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n462_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT93), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n463_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G228gat), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(G78gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(new_n250_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n358_), .B1(new_n389_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G22gat), .B(G50gat), .Z(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(new_n474_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n466_), .A2(new_n469_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n479_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n441_), .A2(new_n461_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n369_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n371_), .A2(KEYINPUT27), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT27), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n488_), .A2(new_n489_), .B1(new_n490_), .B2(new_n372_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n484_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n492_), .A2(new_n459_), .A3(new_n457_), .A4(new_n482_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n460_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n429_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G120gat), .B(G148gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT5), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G176gat), .B(G204gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  NAND2_X1  g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT64), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G57gat), .B(G64gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT71), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(KEYINPUT11), .B2(new_n505_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n508_), .B(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n243_), .B(new_n511_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n261_), .B1(new_n269_), .B2(new_n245_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n220_), .B1(new_n514_), .B2(new_n266_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n282_), .B1(new_n515_), .B2(new_n244_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n511_), .B1(new_n516_), .B2(new_n243_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n504_), .B1(new_n513_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT72), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT72), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n520_), .B(new_n504_), .C1(new_n513_), .C2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n511_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n272_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(KEYINPUT12), .A3(new_n512_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n272_), .A2(new_n526_), .A3(new_n523_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n504_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n502_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n504_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n512_), .A2(KEYINPUT12), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n517_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n527_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n502_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n521_), .A3(new_n519_), .A4(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(KEYINPUT13), .A3(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT82), .B(G15gat), .ZN(new_n542_));
  INV_X1    g341(.A(G22gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT83), .B(G1gat), .Z(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(G8gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G8gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n544_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n284_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n551_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n275_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT86), .ZN(new_n558_));
  INV_X1    g357(.A(new_n553_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n556_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n554_), .A2(new_n555_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT86), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n552_), .A2(new_n563_), .A3(new_n553_), .A4(new_n556_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G113gat), .B(G141gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT87), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G169gat), .B(G197gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n558_), .A2(new_n562_), .A3(new_n564_), .A4(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n541_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n498_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n554_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n523_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT85), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n578_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n306_), .A2(new_n575_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n592_), .A2(new_n546_), .A3(new_n496_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT38), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT100), .Z(new_n596_));
  INV_X1    g395(.A(new_n302_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n498_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n590_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n574_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n429_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n594_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n596_), .A2(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(new_n601_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G8gat), .B1(new_n605_), .B2(new_n491_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT39), .Z(new_n607_));
  NOR3_X1   g406(.A1(new_n592_), .A2(G8gat), .A3(new_n491_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n605_), .B2(new_n461_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT41), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n592_), .A2(G15gat), .A3(new_n461_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT101), .Z(G1326gat));
  XOR2_X1   g414(.A(new_n485_), .B(KEYINPUT102), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n543_), .B1(new_n601_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT42), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n543_), .A3(new_n617_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1327gat));
  NAND3_X1  g420(.A1(new_n487_), .A2(KEYINPUT103), .A3(new_n497_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623_));
  INV_X1    g422(.A(new_n497_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n486_), .A2(new_n461_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n425_), .B2(new_n440_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n304_), .A2(new_n305_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT43), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT43), .B1(new_n487_), .B2(new_n497_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n306_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n498_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT104), .B1(new_n635_), .B2(new_n629_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(new_n633_), .A3(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n599_), .A2(new_n541_), .A3(new_n573_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT44), .B1(new_n637_), .B2(new_n638_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n640_), .A2(new_n496_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G29gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n575_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n597_), .A2(new_n599_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT105), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n429_), .A2(new_n643_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT106), .Z(new_n652_));
  OAI22_X1  g451(.A1(new_n642_), .A2(new_n643_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(new_n650_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n491_), .A2(G36gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT45), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT45), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n660_), .A3(new_n657_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n659_), .A2(new_n661_), .B1(KEYINPUT108), .B2(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(KEYINPUT108), .ZN(new_n664_));
  INV_X1    g463(.A(new_n641_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n491_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n639_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G36gat), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n663_), .A2(new_n664_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n664_), .B1(new_n663_), .B2(new_n668_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  NOR2_X1   g470(.A1(new_n640_), .A2(new_n641_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n461_), .A2(new_n448_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT109), .B(G43gat), .Z(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n656_), .B2(new_n460_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n674_), .A2(KEYINPUT47), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT47), .B1(new_n674_), .B2(new_n676_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1330gat));
  OR3_X1    g478(.A1(new_n650_), .A2(G50gat), .A3(new_n616_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n672_), .A2(new_n681_), .A3(new_n485_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n672_), .B2(new_n485_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1331gat));
  INV_X1    g484(.A(new_n573_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n590_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n541_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n598_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n496_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n541_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n686_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n498_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n629_), .A3(new_n599_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT111), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n496_), .A2(G57gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n691_), .B1(new_n697_), .B2(new_n698_), .ZN(G1332gat));
  INV_X1    g498(.A(G64gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n689_), .B2(new_n666_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT48), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n696_), .A2(new_n700_), .A3(new_n666_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1333gat));
  OAI21_X1  g503(.A(G71gat), .B1(new_n690_), .B2(new_n461_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT49), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n461_), .A2(G71gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n697_), .B2(new_n707_), .ZN(G1334gat));
  AOI21_X1  g507(.A(new_n472_), .B1(new_n689_), .B2(new_n617_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT50), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n696_), .A2(new_n472_), .A3(new_n617_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n692_), .A2(new_n599_), .A3(new_n686_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n637_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G85gat), .B1(new_n715_), .B2(new_n496_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n694_), .A2(new_n645_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n216_), .A3(new_n429_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1336gat));
  OAI21_X1  g518(.A(G92gat), .B1(new_n715_), .B2(new_n491_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n217_), .A3(new_n666_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1337gat));
  AOI21_X1  g521(.A(new_n249_), .B1(new_n714_), .B2(new_n460_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n461_), .A2(new_n224_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n717_), .B2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g525(.A1(new_n637_), .A2(new_n485_), .A3(new_n713_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT114), .B1(new_n727_), .B2(G106gat), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n728_), .A2(new_n729_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n717_), .A2(new_n250_), .A3(new_n485_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT112), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .A4(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n732_), .A2(new_n731_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(new_n737_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT53), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1339gat));
  NAND2_X1  g542(.A1(new_n692_), .A2(new_n687_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n692_), .A2(new_n687_), .A3(KEYINPUT115), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n629_), .A3(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n746_), .A2(new_n629_), .A3(new_n747_), .A4(new_n749_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n536_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n552_), .A2(new_n559_), .A3(new_n556_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n553_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n569_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n572_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n754_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n525_), .A2(new_n504_), .A3(new_n527_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n534_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n528_), .A2(KEYINPUT117), .A3(KEYINPUT55), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT55), .B(new_n530_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n763_), .A3(new_n766_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n502_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n502_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n759_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT58), .B(new_n759_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n772_), .A2(new_n304_), .A3(new_n305_), .A4(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n573_), .A2(new_n754_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n758_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT118), .B1(new_n537_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n779_), .B(new_n758_), .C1(new_n529_), .C2(new_n536_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT57), .B(new_n302_), .C1(new_n776_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n776_), .A2(new_n781_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n597_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n774_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n590_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n753_), .B1(new_n787_), .B2(KEYINPUT120), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n590_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT59), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n666_), .A2(new_n496_), .A3(new_n494_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n786_), .A2(KEYINPUT119), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n774_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n590_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n753_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n793_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n801_), .B2(new_n792_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802_), .B2(new_n573_), .ZN(new_n803_));
  INV_X1    g602(.A(G113gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n801_), .A2(new_n804_), .A3(new_n686_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1340gat));
  OAI21_X1  g605(.A(G120gat), .B1(new_n802_), .B2(new_n692_), .ZN(new_n807_));
  INV_X1    g606(.A(G120gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n692_), .B2(KEYINPUT60), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n801_), .B(new_n809_), .C1(KEYINPUT60), .C2(new_n808_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1341gat));
  OAI21_X1  g610(.A(G127gat), .B1(new_n802_), .B2(new_n590_), .ZN(new_n812_));
  INV_X1    g611(.A(G127gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n801_), .A2(new_n813_), .A3(new_n599_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1342gat));
  NAND2_X1  g614(.A1(new_n801_), .A2(new_n302_), .ZN(new_n816_));
  INV_X1    g615(.A(G134gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT121), .B(G134gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n306_), .A2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT122), .Z(new_n821_));
  OAI211_X1 g620(.A(new_n794_), .B(new_n821_), .C1(new_n801_), .C2(new_n792_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n818_), .A2(new_n822_), .ZN(G1343gat));
  AOI21_X1  g622(.A(new_n493_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n666_), .A2(new_n496_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n686_), .A3(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n541_), .A3(new_n825_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n825_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n590_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT61), .B(G155gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1346gat));
  OAI21_X1  g632(.A(G162gat), .B1(new_n830_), .B2(new_n629_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n597_), .A2(G162gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n830_), .B2(new_n835_), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n491_), .A2(new_n429_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n460_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT123), .Z(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n617_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n330_), .B1(new_n842_), .B2(new_n686_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(KEYINPUT62), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n686_), .A3(new_n347_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(KEYINPUT62), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(G1348gat));
  AOI21_X1  g646(.A(G176gat), .B1(new_n842_), .B2(new_n541_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n839_), .A2(new_n331_), .A3(new_n692_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT124), .B1(new_n800_), .B2(new_n486_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n851_), .B(new_n485_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT125), .B(new_n849_), .C1(new_n850_), .C2(new_n852_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n848_), .B1(new_n855_), .B2(new_n856_), .ZN(G1349gat));
  NOR2_X1   g656(.A1(new_n590_), .A2(new_n340_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n791_), .A2(new_n840_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT126), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n842_), .A2(new_n861_), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n839_), .A2(new_n590_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n321_), .B2(new_n865_), .ZN(G1350gat));
  INV_X1    g665(.A(KEYINPUT127), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n302_), .A2(new_n341_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n842_), .A2(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n842_), .A2(new_n306_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n867_), .B(new_n869_), .C1(new_n870_), .C2(new_n322_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n869_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n322_), .B1(new_n842_), .B2(new_n306_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT127), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1351gat));
  NAND2_X1  g674(.A1(new_n824_), .A2(new_n837_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n573_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n312_), .ZN(G1352gat));
  INV_X1    g677(.A(new_n876_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G204gat), .B1(new_n879_), .B2(new_n541_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n876_), .A2(new_n692_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n310_), .B2(new_n881_), .ZN(G1353gat));
  XOR2_X1   g681(.A(KEYINPUT63), .B(G211gat), .Z(new_n883_));
  NAND3_X1  g682(.A1(new_n879_), .A2(new_n599_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n876_), .B2(new_n590_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1354gat));
  OR3_X1    g686(.A1(new_n876_), .A2(G218gat), .A3(new_n597_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G218gat), .B1(new_n876_), .B2(new_n629_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1355gat));
endmodule


