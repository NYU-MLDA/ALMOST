//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n782_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203_));
  XOR2_X1   g002(.A(G120gat), .B(G148gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G176gat), .B(G204gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT73), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(KEYINPUT11), .ZN(new_n213_));
  INV_X1    g012(.A(G64gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G57gat), .ZN(new_n215_));
  INV_X1    g014(.A(G57gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G64gat), .ZN(new_n217_));
  AND4_X1   g016(.A1(new_n211_), .A2(new_n215_), .A3(new_n217_), .A4(KEYINPUT11), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT68), .B1(new_n213_), .B2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G71gat), .B(G78gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT11), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT69), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n215_), .A2(new_n217_), .A3(new_n211_), .A4(KEYINPUT11), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n219_), .A2(new_n222_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n222_), .B1(new_n219_), .B2(new_n227_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT6), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n238_), .A2(KEYINPUT6), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n231_), .B(new_n235_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G85gat), .B(G92gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT8), .ZN(new_n244_));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n245_));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(new_n241_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n240_), .A2(new_n248_), .A3(KEYINPUT67), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n240_), .B2(new_n248_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n244_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT10), .B(G99gat), .ZN(new_n252_));
  OAI22_X1  g051(.A1(new_n252_), .A2(G106gat), .B1(new_n237_), .B2(new_n239_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G85gat), .A2(G92gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G85gat), .A2(G92gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n256_), .B2(KEYINPUT9), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT9), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n262_), .B2(KEYINPUT65), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n257_), .B(new_n264_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n230_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n251_), .B(new_n266_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(new_n274_), .A3(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n240_), .A2(new_n248_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n240_), .A2(new_n248_), .A3(KEYINPUT67), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n280_), .A2(new_n244_), .B1(new_n265_), .B2(new_n263_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n222_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n225_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n219_), .A2(new_n222_), .A3(new_n227_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n281_), .A2(KEYINPUT12), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(new_n230_), .B2(new_n267_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n275_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n274_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n273_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n268_), .A2(KEYINPUT12), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n230_), .A2(new_n267_), .A3(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n292_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n275_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT71), .B1(new_n300_), .B2(new_n273_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n203_), .B(new_n210_), .C1(new_n295_), .C2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n293_), .A2(new_n208_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n293_), .A2(new_n294_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(KEYINPUT71), .A3(new_n273_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n203_), .B1(new_n308_), .B2(new_n210_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n305_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n209_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n303_), .B1(new_n312_), .B2(new_n203_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n210_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT74), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT75), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n202_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n310_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(KEYINPUT75), .A3(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT13), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G29gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT78), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G43gat), .B(G50gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT15), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G8gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT82), .ZN(new_n328_));
  INV_X1    g127(.A(G15gat), .ZN(new_n329_));
  INV_X1    g128(.A(G22gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G15gat), .A2(G22gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G1gat), .A2(G8gat), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n331_), .A2(new_n332_), .B1(KEYINPUT14), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n328_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n326_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n325_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n325_), .B(new_n335_), .Z(new_n341_));
  INV_X1    g140(.A(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G113gat), .B(G141gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(G169gat), .B(G197gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n344_), .B(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n321_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT105), .ZN(new_n350_));
  OR2_X1    g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  OR2_X1    g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT92), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n353_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT2), .Z(new_n358_));
  OAI211_X1 g157(.A(new_n351_), .B(new_n352_), .C1(new_n356_), .C2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(KEYINPUT1), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n351_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n352_), .A2(KEYINPUT1), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n353_), .B(new_n357_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT91), .ZN(new_n368_));
  XOR2_X1   g167(.A(G113gat), .B(G120gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n364_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n373_), .B2(new_n366_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G85gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT0), .B(G57gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NOR2_X1   g180(.A1(new_n372_), .A2(new_n376_), .ZN(new_n382_));
  OR4_X1    g181(.A1(new_n350_), .A2(new_n377_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n374_), .A2(new_n376_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n381_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n385_), .B(new_n386_), .C1(new_n376_), .C2(new_n372_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n350_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT88), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT99), .ZN(new_n391_));
  INV_X1    g190(.A(G176gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n390_), .A2(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT23), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(G183gat), .B2(G190gat), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n394_), .B(new_n397_), .C1(new_n391_), .C2(new_n390_), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n395_), .B(KEYINPUT23), .Z(new_n399_));
  NOR2_X1   g198(.A1(G169gat), .A2(G176gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT24), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n402_), .A2(new_n403_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n389_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT26), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT26), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT98), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n398_), .B1(new_n407_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G197gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n417_), .A2(G204gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(G204gat), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT21), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G211gat), .B(G218gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(KEYINPUT94), .B2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(KEYINPUT94), .B2(new_n419_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n420_), .B(new_n421_), .C1(new_n423_), .C2(KEYINPUT21), .ZN(new_n424_));
  INV_X1    g223(.A(new_n421_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(KEYINPUT21), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n416_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n408_), .A2(KEYINPUT86), .A3(G190gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n412_), .B2(KEYINPUT86), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT25), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G183gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT84), .B(G183gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n430_), .B(new_n434_), .C1(new_n431_), .C2(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n404_), .B(new_n437_), .C1(new_n405_), .C2(new_n390_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n396_), .B1(new_n436_), .B2(G190gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT90), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n393_), .A2(KEYINPUT89), .ZN(new_n441_));
  INV_X1    g240(.A(G169gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT22), .ZN(new_n443_));
  AOI21_X1  g242(.A(G176gat), .B1(new_n443_), .B2(KEYINPUT89), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n390_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n396_), .B(new_n446_), .C1(new_n436_), .C2(G190gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n438_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n428_), .B(KEYINPUT20), .C1(new_n427_), .C2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT19), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT100), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n449_), .B2(new_n427_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n452_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n457_), .B(new_n458_), .C1(new_n427_), .C2(new_n416_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G8gat), .B(G36gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G64gat), .B(G92gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT32), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n455_), .A2(new_n459_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n427_), .B1(new_n416_), .B2(KEYINPUT104), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(KEYINPUT104), .B2(new_n416_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n457_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n452_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n452_), .B2(new_n450_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT32), .A3(new_n464_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n383_), .A2(new_n388_), .A3(new_n466_), .A4(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(KEYINPUT102), .A2(KEYINPUT33), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n384_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n384_), .A2(new_n474_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n374_), .A2(new_n376_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT103), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n386_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n475_), .B(new_n476_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n455_), .A2(new_n459_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n464_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n455_), .A2(new_n464_), .A3(new_n459_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n473_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n487_));
  OAI21_X1  g286(.A(new_n427_), .B1(new_n364_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G228gat), .A2(G233gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT93), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n427_), .B(new_n490_), .C1(new_n364_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G78gat), .B(G106gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT96), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n495_), .B(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT97), .B1(new_n495_), .B2(new_n498_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n364_), .A2(new_n493_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G22gat), .B(G50gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT28), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n501_), .B(new_n503_), .ZN(new_n504_));
  OR3_X1    g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n499_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G71gat), .B(G99gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G43gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n449_), .B(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n510_), .B(new_n370_), .Z(new_n511_));
  NAND2_X1  g310(.A1(G227gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(new_n329_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT30), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT31), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n507_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n486_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT27), .B1(new_n483_), .B2(new_n484_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n464_), .B(KEYINPUT106), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n471_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n484_), .A2(KEYINPUT27), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n383_), .A2(new_n388_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n518_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n507_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n505_), .A2(new_n506_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n518_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n526_), .B(new_n527_), .C1(new_n530_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n520_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n349_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n326_), .A2(new_n267_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n281_), .A2(new_n325_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n537_), .B(new_n538_), .C1(KEYINPUT35), .C2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT35), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT77), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n542_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT79), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT36), .Z(new_n550_));
  OR2_X1    g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT80), .B(KEYINPUT36), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT81), .Z(new_n554_));
  NAND2_X1  g353(.A1(new_n545_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n335_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n230_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT16), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT83), .Z(new_n568_));
  AND2_X1   g367(.A1(new_n564_), .A2(new_n565_), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n560_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n557_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n536_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT107), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(G1gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n527_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT108), .B(KEYINPUT38), .Z(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n535_), .A2(new_n556_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n571_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n349_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n527_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT109), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(new_n582_), .A3(new_n587_), .ZN(G1324gat));
  INV_X1    g387(.A(G8gat), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n483_), .A2(new_n484_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n524_), .B1(new_n590_), .B2(KEYINPUT27), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n576_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n584_), .A2(new_n349_), .A3(new_n591_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(G8gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n593_), .A3(G8gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n592_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(G1325gat));
  OAI21_X1  g399(.A(G15gat), .B1(new_n585_), .B2(new_n528_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT41), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n576_), .A2(new_n329_), .A3(new_n518_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1326gat));
  OAI21_X1  g403(.A(G22gat), .B1(new_n585_), .B2(new_n531_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT110), .B(KEYINPUT42), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n576_), .A2(new_n330_), .A3(new_n507_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  NOR3_X1   g408(.A1(new_n536_), .A2(new_n556_), .A3(new_n572_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n611_), .A2(G29gat), .A3(new_n527_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT44), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n556_), .B(KEYINPUT37), .Z(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n535_), .B2(new_n615_), .ZN(new_n616_));
  AOI211_X1 g415(.A(KEYINPUT43), .B(new_n557_), .C1(new_n520_), .C2(new_n534_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n571_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n349_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n613_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n535_), .A2(new_n615_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT43), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n535_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n624_), .A2(KEYINPUT44), .A3(new_n571_), .A4(new_n349_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n620_), .A2(new_n625_), .A3(new_n578_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n626_), .A2(KEYINPUT111), .A3(G29gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT111), .B1(new_n626_), .B2(G29gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n612_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  NAND2_X1  g428(.A1(new_n620_), .A2(new_n625_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G36gat), .B1(new_n630_), .B2(new_n526_), .ZN(new_n631_));
  INV_X1    g430(.A(G36gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n610_), .A2(new_n632_), .A3(new_n591_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n631_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n631_), .A2(KEYINPUT46), .A3(new_n635_), .A4(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  NAND2_X1  g440(.A1(new_n518_), .A2(G43gat), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n611_), .A2(new_n528_), .ZN(new_n643_));
  OAI22_X1  g442(.A1(new_n630_), .A2(new_n642_), .B1(G43gat), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g444(.A(G50gat), .B1(new_n630_), .B2(new_n531_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n531_), .A2(G50gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT113), .Z(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n611_), .B2(new_n648_), .ZN(G1331gat));
  INV_X1    g448(.A(new_n348_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n321_), .ZN(new_n651_));
  NOR4_X1   g450(.A1(new_n583_), .A2(new_n571_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(G57gat), .A3(new_n578_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT115), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n535_), .A2(new_n348_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n655_), .A2(new_n573_), .A3(new_n651_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n578_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT114), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(new_n658_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n654_), .A2(new_n659_), .A3(new_n660_), .ZN(G1332gat));
  AOI21_X1  g460(.A(new_n214_), .B1(new_n652_), .B2(new_n591_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT48), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(new_n214_), .A3(new_n591_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1333gat));
  INV_X1    g464(.A(G71gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n652_), .B2(new_n518_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT49), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n656_), .A2(new_n666_), .A3(new_n518_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1334gat));
  INV_X1    g469(.A(G78gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n652_), .B2(new_n507_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT50), .Z(new_n673_));
  NAND3_X1  g472(.A1(new_n656_), .A2(new_n671_), .A3(new_n507_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1335gat));
  NOR2_X1   g474(.A1(new_n572_), .A2(new_n650_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n624_), .A2(new_n321_), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G85gat), .B1(new_n677_), .B2(new_n527_), .ZN(new_n678_));
  NOR4_X1   g477(.A1(new_n655_), .A2(new_n556_), .A3(new_n572_), .A4(new_n651_), .ZN(new_n679_));
  INV_X1    g478(.A(G85gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n578_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1336gat));
  OAI21_X1  g481(.A(G92gat), .B1(new_n677_), .B2(new_n526_), .ZN(new_n683_));
  INV_X1    g482(.A(G92gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n679_), .A2(new_n684_), .A3(new_n591_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT116), .Z(G1337gat));
  NOR2_X1   g486(.A1(new_n528_), .A2(new_n252_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT118), .B1(new_n679_), .B2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n624_), .A2(new_n321_), .A3(new_n518_), .A4(new_n676_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT117), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(G99gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n690_), .B2(G99gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g494(.A1(new_n679_), .A2(new_n234_), .A3(new_n507_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n624_), .A2(new_n321_), .A3(new_n507_), .A4(new_n676_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(new_n698_), .A3(G106gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G106gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g501(.A(new_n344_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n347_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n336_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n347_), .B1(new_n341_), .B2(new_n339_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT55), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n300_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n298_), .A2(new_n269_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n272_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n300_), .A2(new_n710_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n210_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n303_), .B1(new_n716_), .B2(KEYINPUT56), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT120), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n348_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT56), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n715_), .A2(KEYINPUT120), .A3(new_n720_), .A4(new_n210_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n717_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n556_), .B1(new_n709_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT57), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT57), .B(new_n556_), .C1(new_n709_), .C2(new_n722_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n716_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n708_), .B1(new_n727_), .B2(new_n720_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n717_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT58), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(KEYINPUT58), .A3(new_n717_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n615_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n725_), .A2(new_n726_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n571_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT54), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n571_), .A2(new_n650_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n317_), .A2(new_n320_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT119), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n317_), .A2(new_n740_), .A3(new_n320_), .A4(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n736_), .B1(new_n742_), .B2(new_n557_), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT54), .B(new_n615_), .C1(new_n739_), .C2(new_n741_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n735_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n591_), .A2(new_n527_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n533_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(KEYINPUT59), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n743_), .A2(new_n744_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT121), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n572_), .B1(new_n734_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n751_), .B2(new_n734_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n747_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT59), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n749_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G113gat), .B1(new_n756_), .B2(new_n348_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n753_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n747_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OR3_X1    g559(.A1(new_n760_), .A2(G113gat), .A3(new_n348_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n761_), .ZN(G1340gat));
  OAI21_X1  g561(.A(G120gat), .B1(new_n756_), .B2(new_n651_), .ZN(new_n763_));
  INV_X1    g562(.A(G120gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n651_), .B2(KEYINPUT60), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n754_), .B(new_n765_), .C1(KEYINPUT60), .C2(new_n764_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(G1341gat));
  OAI21_X1  g566(.A(G127gat), .B1(new_n756_), .B2(new_n571_), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n760_), .A2(G127gat), .A3(new_n571_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1342gat));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n556_), .B(new_n747_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G134gat), .ZN(new_n773_));
  INV_X1    g572(.A(G134gat), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT122), .B(new_n774_), .C1(new_n760_), .C2(new_n556_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n760_), .A2(KEYINPUT59), .B1(new_n745_), .B2(new_n748_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n557_), .A2(new_n774_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n773_), .A2(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(G1343gat));
  AOI21_X1  g577(.A(new_n529_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n650_), .A3(new_n746_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n321_), .A3(new_n746_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g582(.A1(new_n779_), .A2(new_n572_), .A3(new_n746_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT61), .B(G155gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(G1346gat));
  AND2_X1   g585(.A1(new_n779_), .A2(new_n746_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n615_), .A2(G162gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT123), .ZN(new_n789_));
  INV_X1    g588(.A(new_n556_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n779_), .A2(new_n790_), .A3(new_n746_), .ZN(new_n791_));
  INV_X1    g590(.A(G162gat), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n787_), .A2(new_n789_), .B1(new_n791_), .B2(new_n792_), .ZN(G1347gat));
  NAND3_X1  g592(.A1(new_n591_), .A2(new_n527_), .A3(new_n518_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT124), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n526_), .A2(new_n578_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT124), .A3(new_n518_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n507_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n745_), .A2(new_n650_), .A3(new_n393_), .A4(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT62), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n799_), .A2(KEYINPUT125), .A3(new_n650_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT125), .B1(new_n799_), .B2(new_n650_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n507_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n745_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n803_), .B1(new_n807_), .B2(G169gat), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT62), .B(new_n442_), .C1(new_n745_), .C2(new_n806_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n802_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT126), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT126), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n802_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1348gat));
  INV_X1    g613(.A(new_n745_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n801_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n392_), .A3(new_n321_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n507_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n819_), .A2(new_n321_), .A3(new_n799_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n820_), .B2(new_n392_), .ZN(G1349gat));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n572_), .A3(new_n799_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n571_), .A2(new_n414_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n822_), .A2(new_n435_), .B1(new_n817_), .B2(new_n823_), .ZN(G1350gat));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n790_), .A3(new_n413_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n815_), .A2(new_n557_), .A3(new_n816_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n410_), .B2(new_n826_), .ZN(G1351gat));
  NAND3_X1  g626(.A1(new_n779_), .A2(new_n650_), .A3(new_n797_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n417_), .A2(KEYINPUT127), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT127), .B(G197gat), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n828_), .B2(new_n831_), .ZN(G1352gat));
  NAND3_X1  g631(.A1(new_n779_), .A2(new_n321_), .A3(new_n797_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g633(.A1(new_n779_), .A2(new_n572_), .A3(new_n797_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT63), .B(G211gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n835_), .B2(new_n838_), .ZN(G1354gat));
  NAND2_X1  g638(.A1(new_n779_), .A2(new_n797_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G218gat), .B1(new_n840_), .B2(new_n557_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n556_), .A2(G218gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n840_), .B2(new_n842_), .ZN(G1355gat));
endmodule


