//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n204_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(new_n212_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G229gat), .A2(G233gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n214_), .B(new_n212_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G113gat), .B(G141gat), .Z(new_n222_));
  XNOR2_X1  g021(.A(G169gat), .B(G197gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G85gat), .B(G92gat), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT9), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT9), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G85gat), .A3(G92gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT6), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT7), .ZN(new_n239_));
  INV_X1    g038(.A(G99gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n227_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n239_), .A2(new_n240_), .A3(new_n227_), .A4(KEYINPUT64), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n234_), .A2(new_n238_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n237_), .B1(new_n245_), .B2(new_n229_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n236_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n252_));
  XOR2_X1   g051(.A(G71gat), .B(G78gat), .Z(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(KEYINPUT66), .A3(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n245_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n235_), .B1(new_n258_), .B2(new_n246_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n256_), .B(new_n235_), .C1(new_n258_), .C2(new_n246_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n257_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT67), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT67), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n259_), .A2(new_n260_), .B1(new_n271_), .B2(KEYINPUT12), .ZN(new_n272_));
  INV_X1    g071(.A(new_n261_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n262_), .A2(new_n266_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n269_), .A2(new_n270_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G176gat), .B(G204gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n271_), .A2(KEYINPUT12), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n261_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n259_), .A2(new_n260_), .A3(new_n274_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n276_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n270_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n268_), .A2(KEYINPUT67), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n281_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n283_), .A2(new_n291_), .A3(KEYINPUT13), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(KEYINPUT69), .A3(new_n294_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n225_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G183gat), .ZN(new_n303_));
  INV_X1    g102(.A(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308_));
  INV_X1    g107(.A(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT24), .A3(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n303_), .B2(KEYINPUT78), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(KEYINPUT79), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n325_), .A2(new_n327_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n314_), .B1(new_n323_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT80), .B(G43gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n333_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(G15gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT30), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n337_), .B(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT83), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(KEYINPUT83), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G127gat), .B(G134gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n346_), .A2(new_n347_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n348_), .B1(new_n351_), .B2(new_n345_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT82), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n343_), .A2(new_n344_), .A3(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n354_), .A2(new_n344_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(G211gat), .B(G218gat), .Z(new_n360_));
  OR2_X1    g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n360_), .A2(KEYINPUT21), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(KEYINPUT21), .A3(new_n362_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT21), .ZN(new_n365_));
  AND2_X1   g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G197gat), .A2(G204gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G211gat), .B(G218gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  INV_X1    g171(.A(G141gat), .ZN(new_n373_));
  INV_X1    g172(.A(G148gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT84), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(G155gat), .A3(G162gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n380_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n384_), .A3(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n389_), .A2(new_n386_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT85), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n385_), .B2(KEYINPUT1), .ZN(new_n392_));
  AOI211_X1 g191(.A(KEYINPUT85), .B(new_n388_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n373_), .A2(new_n374_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n387_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n371_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G78gat), .ZN(new_n401_));
  INV_X1    g200(.A(G78gat), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n402_), .B(new_n371_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n401_), .A2(G106gat), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(G106gat), .B1(new_n401_), .B2(new_n403_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n359_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n387_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n389_), .A2(new_n386_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n385_), .A2(KEYINPUT1), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT85), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n385_), .A2(new_n391_), .A3(KEYINPUT1), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n397_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n407_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT28), .B1(new_n414_), .B2(KEYINPUT29), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n371_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(KEYINPUT86), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT28), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n398_), .A2(new_n419_), .A3(new_n399_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n415_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n414_), .A2(KEYINPUT29), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n402_), .B1(new_n424_), .B2(new_n371_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n403_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n227_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n401_), .A2(G106gat), .A3(new_n403_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n359_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n406_), .A2(new_n423_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n423_), .B1(new_n406_), .B2(new_n430_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n352_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n414_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n351_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n398_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(KEYINPUT4), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n414_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G85gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT96), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n398_), .A2(new_n352_), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n351_), .B(new_n387_), .C1(new_n394_), .C2(new_n397_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n441_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n442_), .A2(new_n440_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n444_), .B(new_n450_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n453_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n450_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(KEYINPUT97), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n460_), .A2(new_n461_), .ZN(new_n465_));
  AOI211_X1 g264(.A(new_n453_), .B(new_n450_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n433_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G64gat), .B(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT19), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n477_), .B(KEYINPUT87), .Z(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT88), .B(KEYINPUT20), .C1(new_n333_), .C2(new_n371_), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT25), .B(G183gat), .Z(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT26), .B(G190gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n318_), .A2(new_n319_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n480_), .A2(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n485_));
  OAI21_X1  g284(.A(new_n317_), .B1(new_n485_), .B2(new_n318_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n314_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n371_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n325_), .A2(new_n327_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n330_), .A2(new_n331_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n321_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n320_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n494_), .A2(new_n370_), .A3(new_n363_), .A4(new_n314_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT88), .B1(new_n495_), .B2(KEYINPUT20), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n475_), .B(new_n478_), .C1(new_n489_), .C2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n487_), .A2(new_n371_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n477_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n333_), .A2(new_n371_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n498_), .A2(KEYINPUT20), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n371_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(new_n488_), .A3(new_n479_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n475_), .B1(new_n506_), .B2(new_n478_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n474_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n478_), .B1(new_n489_), .B2(new_n496_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT90), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n510_), .A2(new_n473_), .A3(new_n501_), .A4(new_n497_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(KEYINPUT92), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT27), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n502_), .A2(new_n507_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n473_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n506_), .A2(new_n478_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n498_), .A2(KEYINPUT20), .A3(new_n500_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n477_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT27), .B(new_n511_), .C1(new_n521_), .C2(new_n473_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n468_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n512_), .A2(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n435_), .A2(new_n437_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n451_), .B1(new_n526_), .B2(new_n439_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT95), .B(new_n451_), .C1(new_n526_), .C2(new_n439_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT33), .B1(new_n458_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n458_), .A2(new_n533_), .A3(KEYINPUT33), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n525_), .B(new_n532_), .C1(new_n534_), .C2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n473_), .A2(KEYINPUT32), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n538_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n514_), .B2(new_n538_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n459_), .A2(new_n540_), .A3(new_n462_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n433_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n358_), .B1(new_n524_), .B2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n467_), .A2(new_n463_), .A3(new_n357_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n517_), .B(new_n522_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT98), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n467_), .A2(new_n463_), .A3(new_n357_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT98), .B1(new_n549_), .B2(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n299_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n256_), .B(new_n212_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n556_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(KEYINPUT17), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n556_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT77), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n249_), .A2(new_n214_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n205_), .B2(new_n249_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT71), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(KEYINPUT71), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT72), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT73), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n583_), .B(new_n584_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n587_), .A2(new_n589_), .A3(KEYINPUT74), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT74), .B1(new_n587_), .B2(new_n589_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n570_), .A2(new_n579_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n573_), .A2(new_n593_), .A3(new_n575_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n580_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n587_), .B1(new_n580_), .B2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT37), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n587_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n594_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n578_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n587_), .A2(new_n589_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n580_), .A2(new_n594_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n597_), .A2(new_n605_), .A3(KEYINPUT75), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(KEYINPUT75), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n553_), .A2(new_n568_), .A3(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n467_), .A2(new_n463_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n207_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT99), .Z(new_n613_));
  OR2_X1    g412(.A1(new_n613_), .A2(KEYINPUT38), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(KEYINPUT38), .ZN(new_n615_));
  INV_X1    g414(.A(new_n225_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n298_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT69), .B1(new_n293_), .B2(new_n294_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n566_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n601_), .A2(new_n604_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n552_), .A2(KEYINPUT100), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT100), .B1(new_n552_), .B2(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n610_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(new_n615_), .A3(new_n625_), .ZN(G1324gat));
  NAND3_X1  g425(.A1(new_n609_), .A2(new_n208_), .A3(new_n523_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n628_));
  INV_X1    g427(.A(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n523_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n630_), .B2(G8gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT39), .B(new_n208_), .C1(new_n629_), .C2(new_n523_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n627_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n633_), .B(new_n635_), .ZN(G1325gat));
  NAND3_X1  g435(.A1(new_n609_), .A2(new_n339_), .A3(new_n357_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n357_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(new_n638_), .B2(G15gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n609_), .A2(new_n642_), .A3(new_n433_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n629_), .A2(new_n433_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G22gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT103), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n647_), .A3(G22gat), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n649_));
  AND3_X1   g448(.A1(new_n646_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n643_), .B1(new_n650_), .B2(new_n651_), .ZN(G1327gat));
  NOR3_X1   g451(.A1(new_n553_), .A2(new_n567_), .A3(new_n621_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n611_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n547_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n549_), .A2(new_n545_), .A3(KEYINPUT98), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n523_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n610_), .A2(new_n433_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n525_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n532_), .B1(new_n536_), .B2(new_n534_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n541_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n433_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n357_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n655_), .B(new_n608_), .C1(new_n658_), .C2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n552_), .A2(KEYINPUT104), .A3(new_n655_), .A4(new_n608_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n660_), .A2(new_n665_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n671_), .A2(new_n358_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n606_), .A2(new_n607_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n669_), .A2(new_n670_), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n619_), .A2(new_n567_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT44), .B1(new_n675_), .B2(new_n676_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n611_), .A2(G29gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n654_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  NOR2_X1   g480(.A1(new_n619_), .A2(new_n672_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n621_), .A2(new_n567_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n523_), .B(KEYINPUT105), .Z(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .A4(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n299_), .A2(new_n552_), .A3(new_n684_), .A4(new_n686_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT106), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n687_), .A2(new_n689_), .A3(KEYINPUT45), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT45), .B1(new_n687_), .B2(new_n689_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n677_), .A2(new_n678_), .A3(new_n659_), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n696_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n675_), .A2(new_n676_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n676_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n523_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n706_), .A2(new_n697_), .A3(new_n698_), .A4(new_n692_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n700_), .A2(new_n707_), .ZN(G1329gat));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n358_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n679_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n703_), .A2(new_n704_), .A3(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n653_), .A2(new_n357_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n710_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT47), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n712_), .A2(new_n714_), .A3(new_n719_), .A4(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1330gat));
  AOI21_X1  g520(.A(G50gat), .B1(new_n653_), .B2(new_n433_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n433_), .A2(G50gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n679_), .B2(new_n723_), .ZN(G1331gat));
  INV_X1    g523(.A(G57gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n297_), .A2(new_n298_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n672_), .A3(new_n616_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n608_), .A2(new_n568_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n725_), .B(new_n611_), .C1(new_n729_), .C2(KEYINPUT109), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(KEYINPUT109), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n622_), .A2(new_n623_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n726_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n568_), .A2(new_n616_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n732_), .A2(new_n610_), .A3(new_n735_), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n730_), .A2(new_n731_), .B1(new_n736_), .B2(new_n725_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n732_), .A2(new_n735_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n685_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT48), .Z(new_n743_));
  INV_X1    g542(.A(new_n729_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n739_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n740_), .B2(new_n357_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n744_), .A2(new_n747_), .A3(new_n357_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  AOI21_X1  g550(.A(new_n402_), .B1(new_n740_), .B2(new_n433_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n744_), .A2(new_n402_), .A3(new_n433_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NAND2_X1  g554(.A1(new_n727_), .A2(new_n684_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT111), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n611_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n675_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n726_), .A2(new_n567_), .A3(new_n616_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n611_), .A2(G85gat), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT112), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n758_), .B1(new_n762_), .B2(new_n764_), .ZN(G1336gat));
  INV_X1    g564(.A(G92gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n766_), .A3(new_n523_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n759_), .A2(new_n685_), .A3(new_n761_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(new_n768_), .ZN(G1337gat));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n357_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G99gat), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n357_), .A2(new_n226_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT113), .B1(new_n757_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n757_), .A2(new_n227_), .A3(new_n433_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n675_), .A2(new_n433_), .A3(new_n760_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(G106gat), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n777_), .A3(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(new_n295_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT54), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n673_), .A2(new_n783_), .A3(new_n734_), .A4(new_n785_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n734_), .A2(new_n294_), .A3(new_n293_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n608_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n287_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT115), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n287_), .A2(new_n794_), .A3(new_n791_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n285_), .A2(new_n286_), .A3(new_n257_), .A4(new_n264_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n267_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n793_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n275_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n276_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n287_), .B2(new_n791_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n282_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n217_), .A2(new_n220_), .A3(new_n224_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n213_), .A2(new_n215_), .A3(new_n219_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n224_), .B1(new_n218_), .B2(new_n216_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n283_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n804_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n813_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n608_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n225_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n792_), .A2(KEYINPUT115), .B1(new_n267_), .B2(new_n796_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n802_), .A3(new_n795_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT117), .B1(new_n820_), .B2(new_n281_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n818_), .B1(new_n821_), .B2(KEYINPUT56), .ZN(new_n822_));
  AOI211_X1 g621(.A(KEYINPUT117), .B(new_n804_), .C1(new_n820_), .C2(new_n281_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n817_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n804_), .B1(new_n803_), .B2(KEYINPUT117), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(KEYINPUT56), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(KEYINPUT118), .A4(new_n818_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n283_), .A2(new_n291_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n824_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n621_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n830_), .B2(new_n621_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n816_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n790_), .B1(new_n835_), .B2(new_n567_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n610_), .A2(new_n358_), .A3(new_n545_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n790_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n834_), .B2(new_n566_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n838_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n616_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G113gat), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n566_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n830_), .A2(new_n621_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT57), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n830_), .A2(new_n831_), .A3(new_n621_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n848_), .B1(new_n852_), .B2(new_n816_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT119), .B(new_n838_), .C1(new_n853_), .C2(new_n840_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n225_), .A2(G113gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n845_), .A2(new_n856_), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n839_), .A2(new_n733_), .A3(new_n843_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G120gat), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(G120gat), .B1(new_n733_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n860_), .B2(G120gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n847_), .A2(new_n854_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n863_), .ZN(G1341gat));
  AND4_X1   g663(.A1(G127gat), .A2(new_n839_), .A3(new_n848_), .A4(new_n843_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n847_), .A2(new_n854_), .A3(new_n567_), .ZN(new_n866_));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n866_), .A2(new_n870_), .A3(new_n867_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n865_), .B1(new_n869_), .B2(new_n871_), .ZN(G1342gat));
  AND4_X1   g671(.A1(G134gat), .A2(new_n839_), .A3(new_n608_), .A4(new_n843_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n621_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n847_), .A2(new_n854_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(G134gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT121), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n875_), .A2(new_n879_), .A3(new_n876_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n873_), .B1(new_n878_), .B2(new_n880_), .ZN(G1343gat));
  NAND4_X1  g680(.A1(new_n685_), .A2(new_n433_), .A3(new_n611_), .A4(new_n358_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n841_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n616_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(G141gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n733_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n567_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT123), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n883_), .A2(new_n891_), .A3(new_n567_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n883_), .A2(new_n897_), .A3(new_n874_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n841_), .A2(new_n673_), .A3(new_n882_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n685_), .A2(new_n549_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n433_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n836_), .A2(new_n308_), .A3(new_n616_), .A4(new_n903_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n836_), .A2(new_n616_), .A3(new_n905_), .A4(new_n903_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G169gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(new_n311_), .B2(new_n907_), .ZN(G1348gat));
  AND2_X1   g710(.A1(new_n836_), .A2(new_n903_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G176gat), .B1(new_n912_), .B2(new_n733_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n841_), .A2(new_n433_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n726_), .A2(new_n902_), .A3(new_n309_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n567_), .A3(new_n901_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n848_), .A2(new_n480_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n303_), .A2(new_n917_), .B1(new_n912_), .B2(new_n918_), .ZN(G1350gat));
  INV_X1    g718(.A(new_n481_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n912_), .A2(new_n874_), .A3(new_n920_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n912_), .A2(new_n608_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n304_), .ZN(G1351gat));
  NOR2_X1   g722(.A1(new_n468_), .A2(new_n357_), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT125), .Z(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n741_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n841_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n616_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n733_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n848_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AND2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n932_), .B2(new_n933_), .ZN(G1354gat));
  NAND2_X1  g735(.A1(new_n608_), .A2(G218gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT126), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n927_), .A2(new_n938_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n841_), .A2(new_n621_), .A3(new_n926_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


