//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n206_), .A2(new_n210_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n214_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AOI211_X1 g021(.A(KEYINPUT8), .B(new_n218_), .C1(new_n222_), .C2(new_n206_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n208_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n204_), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n219_), .B(new_n227_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n218_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n224_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n223_), .A2(new_n232_), .A3(KEYINPUT65), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n203_), .A2(new_n205_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n219_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n231_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT8), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(new_n224_), .A3(new_n231_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n217_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G64gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G78gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n246_));
  INV_X1    g045(.A(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n243_), .A2(KEYINPUT11), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n245_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT12), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(new_n242_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n217_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT65), .B1(new_n223_), .B2(new_n232_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n238_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n258_), .B2(new_n252_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT64), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n217_), .B1(new_n223_), .B2(new_n232_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT12), .B1(new_n262_), .B2(new_n251_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n250_), .B(new_n217_), .C1(new_n223_), .C2(new_n232_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n254_), .A2(new_n259_), .A3(new_n261_), .A4(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n261_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n255_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(new_n250_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n270_), .B2(new_n265_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G176gat), .B(G204gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n267_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT13), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G229gat), .A2(G233gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G29gat), .B(G36gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G1gat), .B(G8gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(G22gat), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G22gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT14), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(G1gat), .B2(G8gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n292_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  AOI211_X1 g103(.A(new_n302_), .B(new_n291_), .C1(new_n295_), .C2(new_n299_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n290_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n297_), .A2(new_n298_), .A3(new_n296_), .ZN(new_n307_));
  AOI21_X1  g106(.A(G22gat), .B1(new_n293_), .B2(new_n294_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n291_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n292_), .A3(new_n303_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n285_), .A2(new_n286_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n287_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n306_), .A2(new_n314_), .A3(KEYINPUT77), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT77), .B1(new_n306_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n284_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT15), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n312_), .A2(KEYINPUT15), .A3(new_n287_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n319_), .B(new_n320_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(new_n283_), .A3(new_n314_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G113gat), .B(G141gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT78), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G169gat), .B(G197gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT79), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n317_), .A2(new_n330_), .A3(new_n322_), .A4(new_n327_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n317_), .A2(new_n322_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n335_), .A2(KEYINPUT80), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(KEYINPUT80), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n282_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342_));
  INV_X1    g141(.A(G43gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT30), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(G15gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n345_), .B(new_n348_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351_));
  INV_X1    g150(.A(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(G190gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n350_), .B(new_n356_), .C1(new_n357_), .C2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G190gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT25), .B1(new_n352_), .B2(KEYINPUT81), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n361_), .B(new_n362_), .C1(new_n363_), .C2(KEYINPUT81), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n354_), .B(new_n355_), .C1(G183gat), .C2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(G169gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372_));
  INV_X1    g171(.A(G169gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT22), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n370_), .B(new_n371_), .C1(new_n372_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n366_), .B(new_n357_), .C1(new_n375_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n365_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n349_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n349_), .A2(new_n380_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT31), .Z(new_n385_));
  XNOR2_X1  g184(.A(G127gat), .B(G134gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT84), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n386_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n388_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n387_), .A2(KEYINPUT85), .A3(new_n389_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n385_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n384_), .B(KEYINPUT31), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n397_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G22gat), .B(G50gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT90), .ZN(new_n405_));
  XOR2_X1   g204(.A(G197gat), .B(G204gat), .Z(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT21), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G211gat), .B(G218gat), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n406_), .A2(KEYINPUT21), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n407_), .A2(new_n409_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n410_), .A2(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G141gat), .A2(G148gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT3), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G141gat), .A2(G148gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT2), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(KEYINPUT1), .B2(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(KEYINPUT1), .B2(new_n422_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n415_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(new_n417_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n419_), .A2(new_n423_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n405_), .B1(new_n414_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n404_), .A2(KEYINPUT90), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n405_), .B(new_n432_), .C1(new_n414_), .C2(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT88), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n403_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n403_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(KEYINPUT88), .A3(new_n442_), .A4(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n428_), .A2(new_n429_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n443_), .A3(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G8gat), .B(G36gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n410_), .A2(new_n411_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n413_), .A2(new_n412_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n459_), .B1(new_n462_), .B2(new_n380_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT93), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G226gat), .A2(G233gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n366_), .A2(KEYINPUT92), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT92), .B1(new_n352_), .B2(new_n353_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n354_), .A2(new_n470_), .A3(new_n355_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n374_), .A2(new_n368_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n377_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n469_), .A2(new_n471_), .A3(new_n357_), .A4(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT25), .B(G183gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n361_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n360_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n414_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .A4(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n463_), .A2(new_n468_), .A3(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT93), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n365_), .A2(new_n379_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n459_), .B1(new_n482_), .B2(new_n414_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n474_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n462_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n468_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n458_), .B(new_n479_), .C1(new_n481_), .C2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT95), .ZN(new_n488_));
  INV_X1    g287(.A(new_n485_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT20), .B1(new_n462_), .B2(new_n380_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n467_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT93), .A3(new_n480_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT95), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n458_), .A4(new_n479_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n479_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n457_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n488_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT96), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n428_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT97), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n390_), .A2(new_n393_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n428_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT97), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n501_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT99), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT98), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n501_), .B(KEYINPUT99), .C1(new_n499_), .C2(new_n504_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n505_), .A2(KEYINPUT4), .ZN(new_n512_));
  INV_X1    g311(.A(new_n509_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G1gat), .B(G29gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(G85gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT0), .B(G57gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n511_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT33), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n513_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n505_), .A2(new_n509_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n488_), .A2(new_n496_), .A3(new_n528_), .A4(new_n494_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT33), .B(new_n520_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n498_), .A2(new_n527_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n524_), .A2(new_n520_), .A3(new_n525_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n526_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n457_), .A2(KEYINPUT32), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n495_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n483_), .A2(new_n468_), .A3(new_n485_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n463_), .A2(new_n478_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n468_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(KEYINPUT32), .A3(new_n457_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n452_), .B1(new_n531_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT27), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n497_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n538_), .B2(new_n458_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n496_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n449_), .A2(new_n532_), .A3(new_n526_), .A4(new_n450_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n402_), .B1(new_n541_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n402_), .A2(new_n533_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n546_), .A2(new_n452_), .A3(KEYINPUT100), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT100), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n497_), .A2(new_n542_), .B1(new_n496_), .B2(new_n544_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n553_), .B2(new_n451_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n341_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT67), .B(KEYINPUT34), .Z(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n269_), .A2(new_n313_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n319_), .A2(new_n320_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n258_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(new_n558_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT36), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT69), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n571_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n575_), .A3(new_n567_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n557_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n568_), .B(KEYINPUT70), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n572_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n568_), .A2(KEYINPUT70), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n580_), .B(new_n572_), .C1(new_n583_), .C2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n578_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n579_), .B1(new_n588_), .B2(new_n557_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT74), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT76), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT17), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n310_), .A2(new_n311_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n250_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n601_), .A2(new_n595_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n589_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n556_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT101), .ZN(new_n608_));
  INV_X1    g407(.A(G1gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n533_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n588_), .A2(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n556_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n533_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(G8gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n608_), .A2(new_n619_), .A3(new_n546_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G8gat), .B1(new_n615_), .B2(new_n553_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(KEYINPUT102), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(KEYINPUT102), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n622_), .A2(new_n623_), .A3(KEYINPUT39), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n620_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n620_), .B(new_n629_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1325gat));
  INV_X1    g432(.A(new_n402_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n608_), .A2(new_n347_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G15gat), .B1(new_n615_), .B2(new_n402_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT41), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(KEYINPUT41), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(new_n637_), .A3(new_n638_), .ZN(G1326gat));
  OR2_X1    g438(.A1(new_n452_), .A2(KEYINPUT104), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n452_), .A2(KEYINPUT104), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G22gat), .B1(new_n615_), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT42), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n608_), .A2(new_n296_), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n605_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n341_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n589_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n589_), .B2(KEYINPUT105), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n650_), .B(new_n652_), .C1(new_n549_), .C2(new_n555_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n652_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n549_), .A2(new_n555_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n589_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n649_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT44), .B(new_n649_), .C1(new_n653_), .C2(new_n656_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n533_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G29gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n588_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n648_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n556_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n616_), .A2(G29gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT106), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n668_), .ZN(G1328gat));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n670_), .A3(new_n546_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n659_), .A2(new_n546_), .A3(new_n660_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT107), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n659_), .A2(new_n676_), .A3(new_n546_), .A4(new_n660_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n673_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT46), .B(new_n673_), .C1(new_n675_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n665_), .A2(new_n343_), .A3(new_n634_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n659_), .A2(new_n634_), .A3(new_n660_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n343_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1330gat));
  INV_X1    g487(.A(G50gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n665_), .A2(new_n689_), .A3(new_n642_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n659_), .A2(KEYINPUT109), .A3(new_n452_), .A4(new_n660_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(G50gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n659_), .A2(new_n452_), .A3(new_n660_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT110), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  AND4_X1   g495(.A1(KEYINPUT110), .A2(new_n695_), .A3(G50gat), .A4(new_n691_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n690_), .B1(new_n696_), .B2(new_n697_), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n281_), .A2(new_n338_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n655_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n614_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n616_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n700_), .A2(new_n606_), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n533_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(new_n546_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n701_), .A2(new_n546_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G64gat), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT48), .B(new_n708_), .C1(new_n701_), .C2(new_n546_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT111), .Z(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n701_), .B2(new_n634_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT49), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n704_), .A2(new_n716_), .A3(new_n634_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n701_), .B2(new_n642_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT50), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n704_), .A2(new_n721_), .A3(new_n642_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1335gat));
  NOR2_X1   g524(.A1(new_n653_), .A2(new_n656_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n699_), .A2(new_n605_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT112), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n727_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n730_), .B(new_n731_), .C1(new_n653_), .C2(new_n656_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n616_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n700_), .A2(new_n664_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n211_), .A3(new_n533_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  OAI21_X1  g537(.A(G92gat), .B1(new_n734_), .B2(new_n553_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n212_), .A3(new_n546_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  XNOR2_X1  g540(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n402_), .B1(new_n728_), .B2(new_n732_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n743_), .A2(new_n226_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n634_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT113), .B1(new_n736_), .B2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n742_), .C1(new_n743_), .C2(new_n226_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n736_), .A2(new_n208_), .A3(new_n452_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n452_), .B(new_n730_), .C1(new_n653_), .C2(new_n656_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g556(.A1(new_n551_), .A2(new_n554_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n634_), .A2(new_n533_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(KEYINPUT59), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT77), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n290_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n313_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n306_), .A2(new_n314_), .A3(KEYINPUT77), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n284_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n321_), .A2(new_n284_), .A3(new_n314_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n326_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT117), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n283_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n770_), .A2(new_n326_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n763_), .B1(new_n332_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n332_), .A2(new_n763_), .A3(new_n777_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n278_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n254_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n268_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT115), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n785_), .A3(new_n268_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n267_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n242_), .B1(new_n241_), .B2(new_n253_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n264_), .B1(new_n270_), .B2(KEYINPUT12), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT55), .A3(new_n261_), .A4(new_n254_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n784_), .A2(new_n786_), .A3(new_n788_), .A4(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n275_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n781_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT120), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n781_), .B(new_n800_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n589_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI221_X4 g604(.A(KEYINPUT118), .B1(new_n772_), .B2(new_n776_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n277_), .B1(new_n806_), .B2(new_n778_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n793_), .A2(new_n275_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n807_), .B1(new_n810_), .B2(new_n794_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n799_), .B1(new_n811_), .B2(new_n800_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n801_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT121), .B(new_n589_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(KEYINPUT58), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n278_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n794_), .B1(new_n796_), .B2(KEYINPUT116), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n782_), .A2(new_n785_), .A3(new_n268_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n785_), .B1(new_n782_), .B2(new_n268_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n267_), .B(KEYINPUT55), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n276_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(KEYINPUT56), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n818_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n280_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n817_), .B(new_n588_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n824_), .B2(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n796_), .A2(KEYINPUT116), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n794_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n834_), .B2(new_n818_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n817_), .B1(new_n835_), .B2(new_n588_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n831_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n648_), .B1(new_n816_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n282_), .A2(new_n338_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n606_), .A2(new_n839_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n840_), .A2(KEYINPUT54), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(KEYINPUT54), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n762_), .B1(new_n838_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n836_), .B1(new_n830_), .B2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT119), .B(new_n817_), .C1(new_n835_), .C2(new_n588_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n814_), .A2(new_n815_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT121), .B1(new_n802_), .B2(new_n589_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n605_), .B1(new_n848_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n843_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n761_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n844_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n339_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n854_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n339_), .A2(G113gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(G1340gat));
  OAI211_X1 g659(.A(new_n282_), .B(new_n844_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G120gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n281_), .A2(KEYINPUT60), .ZN(new_n863_));
  MUX2_X1   g662(.A(new_n863_), .B(KEYINPUT60), .S(G120gat), .Z(new_n864_));
  NAND2_X1  g663(.A1(new_n854_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT122), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n862_), .A2(new_n868_), .A3(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1341gat));
  OAI21_X1  g669(.A(G127gat), .B1(new_n856_), .B2(new_n605_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n605_), .A2(G127gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n858_), .B2(new_n872_), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n856_), .B2(new_n650_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n663_), .A2(G134gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n858_), .B2(new_n875_), .ZN(G1343gat));
  NAND4_X1  g675(.A1(new_n402_), .A2(new_n533_), .A3(new_n452_), .A4(new_n553_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n338_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n282_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n648_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n878_), .A2(new_n886_), .A3(new_n588_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n878_), .A2(new_n589_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n886_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n838_), .A2(new_n843_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n550_), .A2(new_n546_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n642_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n890_), .A2(KEYINPUT123), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n890_), .B2(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n338_), .A3(new_n472_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n890_), .A2(new_n893_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n338_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n900_), .B2(G169gat), .ZN(new_n901_));
  AOI211_X1 g700(.A(KEYINPUT62), .B(new_n373_), .C1(new_n899_), .C2(new_n338_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n897_), .B1(new_n901_), .B2(new_n902_), .ZN(G1348gat));
  NAND2_X1  g702(.A1(new_n896_), .A2(new_n282_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n452_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n891_), .A2(new_n377_), .A3(new_n281_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n377_), .B1(new_n905_), .B2(new_n906_), .ZN(G1349gat));
  NOR2_X1   g706(.A1(new_n605_), .A2(new_n475_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n905_), .A2(new_n546_), .A3(new_n550_), .A4(new_n648_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n896_), .A2(new_n908_), .B1(new_n352_), .B2(new_n909_), .ZN(G1350gat));
  NAND2_X1  g709(.A1(new_n588_), .A2(new_n361_), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT124), .Z(new_n912_));
  NAND2_X1  g711(.A1(new_n896_), .A2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n650_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n353_), .ZN(G1351gat));
  NOR2_X1   g714(.A1(new_n634_), .A2(new_n547_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT125), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n553_), .B(new_n917_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n338_), .ZN(new_n919_));
  INV_X1    g718(.A(G197gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT126), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n918_), .A2(new_n922_), .A3(G197gat), .A4(new_n338_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n920_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n921_), .A2(new_n923_), .A3(new_n924_), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n918_), .A2(new_n282_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g726(.A1(new_n918_), .A2(new_n648_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT63), .B(G211gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n931_));
  INV_X1    g730(.A(G211gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n928_), .A2(KEYINPUT127), .A3(new_n931_), .A4(new_n932_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n930_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n918_), .A2(new_n938_), .A3(new_n588_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n918_), .A2(new_n589_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n938_), .ZN(G1355gat));
endmodule


