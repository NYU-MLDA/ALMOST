//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(G78gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G22gat), .B(G50gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211_));
  INV_X1    g010(.A(G155gat), .ZN(new_n212_));
  INV_X1    g011(.A(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT91), .B1(G155gat), .B2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G141gat), .A2(G148gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT92), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n227_), .A3(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT93), .B(KEYINPUT2), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT94), .B1(new_n230_), .B2(new_n222_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n223_), .A2(KEYINPUT3), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n232_), .A2(new_n234_), .B1(new_n222_), .B2(KEYINPUT2), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT94), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n237_), .A2(KEYINPUT93), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(KEYINPUT93), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n236_), .B(new_n221_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n231_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n216_), .A2(new_n217_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n229_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT28), .B1(new_n244_), .B2(KEYINPUT29), .ZN(new_n245_));
  OR2_X1    g044(.A1(KEYINPUT96), .A2(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(KEYINPUT96), .A2(G204gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(G197gat), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT95), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT95), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G197gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(G204gat), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT21), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n246_), .A2(G197gat), .A3(new_n247_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n252_), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n255_), .B(new_n256_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n255_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(KEYINPUT21), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n226_), .A2(new_n228_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n269_), .A3(new_n267_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n245_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n245_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n210_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n268_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n270_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n269_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n245_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n209_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G85gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G57gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G134gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G113gat), .B(G120gat), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n228_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n227_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n243_), .B(new_n289_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT98), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT89), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n287_), .A2(KEYINPUT89), .A3(new_n288_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n290_), .A2(new_n291_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n243_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT98), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n229_), .A2(new_n301_), .A3(new_n243_), .A4(new_n289_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n293_), .A2(new_n300_), .A3(new_n302_), .A4(KEYINPUT4), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n229_), .A2(new_n243_), .B1(new_n296_), .B2(new_n295_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n293_), .A2(new_n300_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n284_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n284_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n280_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314_));
  AND2_X1   g113(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n316_));
  OAI21_X1  g115(.A(G169gat), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(KEYINPUT86), .B(G169gat), .C1(new_n315_), .C2(new_n316_), .ZN(new_n320_));
  INV_X1    g119(.A(G169gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(G176gat), .B1(new_n321_), .B2(KEYINPUT22), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  OR2_X1    g123(.A1(KEYINPUT84), .A2(KEYINPUT23), .ZN(new_n325_));
  NAND2_X1  g124(.A1(KEYINPUT84), .A2(KEYINPUT23), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n329_), .A2(KEYINPUT23), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n323_), .A2(new_n324_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n324_), .A2(KEYINPUT24), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  MUX2_X1   g136(.A(new_n336_), .B(KEYINPUT24), .S(new_n337_), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  INV_X1    g139(.A(G183gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(KEYINPUT25), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n339_), .B(new_n342_), .C1(new_n343_), .C2(new_n340_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n329_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n328_), .A2(KEYINPUT23), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n338_), .B(new_n344_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n335_), .A2(new_n261_), .A3(new_n347_), .A4(new_n264_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n261_), .A2(new_n264_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n339_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n338_), .A2(new_n330_), .A3(new_n333_), .A4(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n332_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n324_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n348_), .B(KEYINPUT20), .C1(new_n349_), .C2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n349_), .B2(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n335_), .A2(new_n347_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n365_), .B2(new_n265_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n359_), .A2(new_n362_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G8gat), .B(G36gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT18), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n314_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n359_), .A2(new_n362_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n351_), .A2(new_n357_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n265_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT100), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n365_), .A2(new_n265_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n265_), .C2(new_n374_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n373_), .B1(new_n380_), .B2(new_n362_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n372_), .B1(new_n381_), .B2(new_n371_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n359_), .A2(new_n362_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n364_), .A2(new_n366_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n371_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n371_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n383_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n313_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n312_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n386_), .A2(new_n387_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n303_), .B(new_n304_), .C1(KEYINPUT4), .C2(new_n300_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n284_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n304_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n293_), .A2(new_n300_), .A3(new_n302_), .A4(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n308_), .A2(KEYINPUT33), .A3(new_n309_), .A4(new_n284_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n392_), .A2(new_n393_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT101), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n371_), .A2(KEYINPUT32), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n380_), .A2(new_n362_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n401_), .B(new_n403_), .C1(new_n404_), .C2(new_n373_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT101), .B1(new_n381_), .B2(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n367_), .A2(new_n402_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n308_), .A2(new_n309_), .A3(new_n284_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n310_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n400_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n280_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n390_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT87), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT30), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n365_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT88), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G15gat), .B(G43gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n417_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT31), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n297_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n295_), .A2(KEYINPUT31), .A3(new_n296_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n422_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n427_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n202_), .B1(new_n413_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n311_), .A2(new_n312_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n435_), .A2(new_n405_), .A3(new_n408_), .A4(new_n406_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n280_), .B1(new_n436_), .B2(new_n400_), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT103), .B(new_n432_), .C1(new_n437_), .C2(new_n390_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n389_), .A2(KEYINPUT104), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n389_), .A2(KEYINPUT104), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n432_), .A2(new_n280_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT105), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n432_), .A2(new_n435_), .A3(new_n280_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT105), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n446_), .B(new_n447_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n434_), .A2(new_n438_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G15gat), .B(G22gat), .ZN(new_n451_));
  INV_X1    g250(.A(G1gat), .ZN(new_n452_));
  INV_X1    g251(.A(G8gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT14), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G8gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G43gat), .B(G50gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n462_), .A2(KEYINPUT81), .A3(new_n464_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n450_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n461_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n457_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n472_), .A2(new_n462_), .A3(new_n450_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G113gat), .B(G141gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G169gat), .B(G197gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n469_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT82), .B(new_n477_), .C1(new_n469_), .C2(new_n473_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G230gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G71gat), .B(G78gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT11), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n489_));
  INV_X1    g288(.A(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT6), .ZN(new_n495_));
  INV_X1    g294(.A(G85gat), .ZN(new_n496_));
  INV_X1    g295(.A(G92gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT9), .ZN(new_n499_));
  AND2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n498_), .B(new_n499_), .C1(new_n500_), .C2(KEYINPUT64), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n498_), .A2(new_n502_), .A3(KEYINPUT9), .A4(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n206_), .A3(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n495_), .A2(new_n501_), .A3(new_n504_), .A4(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n206_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n494_), .A2(KEYINPUT6), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n510_), .B(new_n513_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT65), .B1(new_n500_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT65), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n498_), .A2(new_n520_), .A3(new_n503_), .ZN(new_n521_));
  AND4_X1   g320(.A1(new_n509_), .A2(new_n517_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n519_), .A2(new_n521_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n509_), .B1(new_n523_), .B2(new_n517_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n493_), .B(new_n508_), .C1(new_n522_), .C2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT66), .ZN(new_n526_));
  INV_X1    g325(.A(new_n508_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n494_), .B(new_n514_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n513_), .A2(new_n510_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n521_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT8), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n509_), .A3(new_n517_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n527_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n493_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n485_), .B1(new_n526_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT12), .B1(new_n534_), .B2(new_n493_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n508_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  INV_X1    g338(.A(new_n493_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n525_), .A2(new_n484_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n525_), .A2(KEYINPUT67), .A3(new_n484_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G120gat), .B(G148gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n536_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT69), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n536_), .A2(new_n555_), .A3(new_n547_), .A4(new_n552_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n536_), .A2(new_n547_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n551_), .B(KEYINPUT68), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT13), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(KEYINPUT13), .A3(new_n560_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n563_), .A2(KEYINPUT70), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT70), .B1(new_n563_), .B2(new_n564_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n483_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n449_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT77), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n534_), .A2(new_n461_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n471_), .A2(new_n538_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(KEYINPUT72), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n574_), .A2(new_n571_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n575_), .B(new_n576_), .C1(KEYINPUT72), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT73), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT36), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n590_));
  NAND4_X1  g389(.A1(new_n580_), .A2(new_n582_), .A3(new_n587_), .A4(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n570_), .B1(new_n592_), .B2(KEYINPUT37), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n589_), .A2(KEYINPUT77), .A3(new_n594_), .A4(new_n591_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n588_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n597_), .B2(KEYINPUT75), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  AOI211_X1 g398(.A(new_n599_), .B(new_n596_), .C1(new_n580_), .C2(new_n582_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT37), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT76), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(KEYINPUT76), .B(KEYINPUT37), .C1(new_n598_), .C2(new_n600_), .ZN(new_n604_));
  AOI221_X4 g403(.A(new_n569_), .B1(new_n593_), .B2(new_n595_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n593_), .A2(new_n595_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT78), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n457_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n540_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT79), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n616_), .B(KEYINPUT17), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT80), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n612_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n609_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n568_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n452_), .A3(new_n435_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n592_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n449_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n567_), .A2(new_n626_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n443_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n630_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n631_), .A2(new_n637_), .A3(new_n638_), .ZN(G1324gat));
  AOI21_X1  g438(.A(new_n453_), .B1(new_n635_), .B2(new_n441_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT39), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n628_), .A2(new_n453_), .A3(new_n441_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(KEYINPUT40), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n635_), .B2(new_n433_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT41), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n628_), .A2(new_n648_), .A3(new_n433_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n635_), .B2(new_n280_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT42), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n628_), .A2(new_n653_), .A3(new_n280_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n434_), .A2(new_n438_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n445_), .A2(new_n448_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n567_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n626_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n592_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT108), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n568_), .A2(new_n666_), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G29gat), .B1(new_n669_), .B2(new_n435_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n567_), .A2(new_n662_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n660_), .A2(new_n673_), .A3(new_n609_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n589_), .A2(new_n599_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n597_), .A2(KEYINPUT75), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n591_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT76), .B1(new_n677_), .B2(KEYINPUT37), .ZN(new_n678_));
  INV_X1    g477(.A(new_n604_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n607_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n569_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n606_), .A2(KEYINPUT78), .A3(new_n607_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n449_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n672_), .B1(new_n674_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT106), .B1(new_n685_), .B2(KEYINPUT44), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n673_), .B1(new_n660_), .B2(new_n609_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n449_), .A2(new_n683_), .A3(KEYINPUT43), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n687_), .B(new_n688_), .C1(new_n691_), .C2(new_n672_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n671_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n685_), .A2(new_n695_), .A3(KEYINPUT44), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n686_), .A2(new_n692_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n435_), .A2(G29gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n670_), .B1(new_n697_), .B2(new_n698_), .ZN(G1328gat));
  XNOR2_X1  g498(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n697_), .B2(new_n441_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n441_), .A2(KEYINPUT109), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n441_), .A2(KEYINPUT109), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n665_), .A2(new_n667_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT110), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n665_), .A2(new_n667_), .A3(new_n709_), .A4(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(KEYINPUT45), .A3(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n700_), .B1(new_n702_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n692_), .A2(new_n686_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n694_), .A2(new_n696_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n441_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G36gat), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT46), .A3(new_n714_), .A4(new_n713_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n721_), .ZN(G1329gat));
  NAND4_X1  g521(.A1(new_n717_), .A2(new_n718_), .A3(G43gat), .A4(new_n433_), .ZN(new_n723_));
  INV_X1    g522(.A(G43gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n668_), .B2(new_n432_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT47), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n728_), .A3(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1330gat));
  AOI21_X1  g529(.A(G50gat), .B1(new_n669_), .B2(new_n280_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n280_), .A2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n697_), .B2(new_n732_), .ZN(G1331gat));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n565_), .A2(new_n566_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n449_), .A2(new_n736_), .A3(new_n483_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(new_n627_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT112), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n435_), .B1(new_n738_), .B2(KEYINPUT112), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n734_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n742_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n483_), .A2(new_n626_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n633_), .A2(new_n735_), .A3(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n443_), .A2(new_n734_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n743_), .A2(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n705_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n746_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n746_), .B2(new_n433_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT49), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n738_), .A2(new_n756_), .A3(new_n433_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1334gat));
  AOI21_X1  g559(.A(new_n204_), .B1(new_n746_), .B2(new_n280_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT50), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n738_), .A2(new_n204_), .A3(new_n280_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n736_), .A2(new_n662_), .A3(new_n483_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n691_), .A2(KEYINPUT115), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n689_), .A2(new_n690_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n443_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n737_), .A2(new_n663_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n496_), .A3(new_n435_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n769_), .B2(new_n705_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n497_), .A3(new_n441_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  OAI211_X1 g576(.A(new_n433_), .B(new_n765_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G99gat), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n772_), .A2(new_n505_), .A3(new_n506_), .A4(new_n433_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT117), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT51), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n779_), .A2(new_n786_), .A3(new_n780_), .A4(new_n781_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n785_), .A3(new_n787_), .ZN(G1338gat));
  NAND3_X1  g587(.A1(new_n772_), .A2(new_n206_), .A3(new_n280_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n765_), .A2(new_n280_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G106gat), .B1(new_n691_), .B2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT52), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT52), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI211_X1 g594(.A(new_n435_), .B(new_n442_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT121), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n467_), .A2(new_n468_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n450_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n450_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n476_), .B1(new_n472_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n478_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT66), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n525_), .B(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n484_), .B1(new_n806_), .B2(new_n542_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n547_), .A2(KEYINPUT55), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n542_), .A2(new_n545_), .A3(new_n809_), .A4(new_n546_), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT118), .B(new_n807_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n810_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n807_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n559_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT56), .B(new_n559_), .C1(new_n811_), .C2(new_n815_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n804_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT58), .B(new_n804_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n609_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n818_), .A2(KEYINPUT119), .A3(new_n820_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n557_), .B(new_n483_), .C1(new_n820_), .C2(KEYINPUT119), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n483_), .A2(new_n557_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n821_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n818_), .A2(KEYINPUT119), .A3(new_n820_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT120), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n803_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n830_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n592_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n826_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n833_), .A2(new_n834_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n836_), .B1(new_n842_), .B2(new_n827_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n632_), .B1(new_n843_), .B2(new_n835_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT57), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n662_), .B1(new_n841_), .B2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n683_), .A2(new_n563_), .A3(new_n564_), .A4(new_n745_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n797_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n609_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n844_), .B2(KEYINPUT57), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n839_), .A2(new_n840_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n626_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n848_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n797_), .C1(new_n851_), .C2(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n854_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n483_), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  INV_X1    g664(.A(new_n797_), .ZN(new_n866_));
  AOI211_X1 g665(.A(new_n862_), .B(new_n866_), .C1(new_n858_), .C2(new_n848_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n867_), .B2(G113gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT122), .B(new_n863_), .C1(new_n850_), .C2(new_n862_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n861_), .A2(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(G1340gat));
  INV_X1    g669(.A(new_n850_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n736_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n871_), .B(new_n873_), .C1(KEYINPUT60), .C2(new_n872_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n736_), .B1(new_n854_), .B2(new_n860_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n872_), .ZN(G1341gat));
  INV_X1    g675(.A(G127gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n871_), .A2(new_n877_), .A3(new_n662_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n626_), .B1(new_n854_), .B2(new_n860_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n877_), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n871_), .A2(new_n881_), .A3(new_n632_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n683_), .B1(new_n854_), .B2(new_n860_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1343gat));
  NOR4_X1   g683(.A1(new_n750_), .A2(new_n443_), .A3(new_n412_), .A4(new_n433_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n859_), .A2(new_n483_), .A3(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n859_), .A2(new_n735_), .A3(new_n885_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n859_), .A2(new_n885_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n626_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT61), .B(G155gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  OAI21_X1  g692(.A(new_n213_), .B1(new_n890_), .B2(new_n592_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n609_), .A2(G162gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT124), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n859_), .A2(new_n885_), .A3(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n894_), .A2(new_n897_), .ZN(G1347gat));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n846_), .A2(new_n849_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n705_), .A2(new_n444_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n862_), .A3(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n903_), .B2(new_n321_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n859_), .A2(new_n901_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT62), .B(G169gat), .C1(new_n905_), .C2(new_n862_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n354_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  NOR2_X1   g707(.A1(new_n900_), .A2(new_n902_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n910_));
  OR2_X1    g709(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n909_), .A2(new_n735_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n905_), .A2(new_n736_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1349gat));
  AOI21_X1  g713(.A(G183gat), .B1(new_n909_), .B2(new_n662_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n905_), .A2(new_n626_), .A3(new_n343_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n909_), .A2(new_n632_), .A3(new_n339_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G190gat), .B1(new_n905_), .B2(new_n683_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n433_), .A2(new_n313_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n750_), .A2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n859_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n862_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n249_), .ZN(G1352gat));
  NAND3_X1  g725(.A1(new_n859_), .A2(new_n735_), .A3(new_n923_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n246_), .A2(new_n247_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n900_), .A2(new_n736_), .A3(new_n922_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n929_), .ZN(new_n932_));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n927_), .A2(G204gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n930_), .B1(new_n933_), .B2(new_n934_), .ZN(G1353gat));
  NOR2_X1   g734(.A1(new_n900_), .A2(new_n922_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n937_));
  INV_X1    g736(.A(G211gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n662_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n937_), .A2(new_n938_), .A3(KEYINPUT127), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n936_), .A2(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n924_), .A2(new_n939_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n943_), .ZN(G1354gat));
  OR3_X1    g745(.A1(new_n924_), .A2(G218gat), .A3(new_n592_), .ZN(new_n947_));
  OAI21_X1  g746(.A(G218gat), .B1(new_n924_), .B2(new_n683_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1355gat));
endmodule


