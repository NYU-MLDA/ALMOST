//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_;
  NAND3_X1  g000(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND4_X1  g003(.A1(KEYINPUT87), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT85), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT3), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n215_), .A2(new_n211_), .A3(new_n212_), .A4(KEYINPUT85), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n206_), .A2(new_n210_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G155gat), .B2(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(G155gat), .ZN(new_n220_));
  INV_X1    g019(.A(G162gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT83), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n219_), .A2(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT1), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(new_n232_), .A3(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(new_n219_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G141gat), .B(G148gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT88), .ZN(new_n239_));
  XOR2_X1   g038(.A(G127gat), .B(G134gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT88), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(new_n237_), .A3(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n238_), .A2(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G225gat), .A2(G233gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT96), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT97), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT97), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n245_), .A2(new_n252_), .A3(new_n246_), .A4(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G85gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n239_), .A2(new_n260_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n261_), .A2(new_n248_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n245_), .A2(KEYINPUT4), .A3(new_n246_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n251_), .A2(new_n253_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n266_), .A2(new_n259_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n239_), .A2(new_n244_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G22gat), .B(G50gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT28), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n270_), .B(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G197gat), .A2(G204gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT21), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278_));
  INV_X1    g077(.A(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n274_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G211gat), .B(G218gat), .Z(new_n283_));
  NAND4_X1  g082(.A1(new_n283_), .A2(KEYINPUT21), .A3(new_n275_), .A4(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT89), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n284_), .A3(KEYINPUT89), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n269_), .B1(new_n228_), .B2(new_n237_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n285_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G78gat), .B(G106gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT90), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n292_), .A2(new_n298_), .A3(new_n295_), .ZN(new_n301_));
  AND4_X1   g100(.A1(KEYINPUT91), .A2(new_n273_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT91), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n304_), .A2(new_n273_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n265_), .B(new_n267_), .C1(new_n302_), .C2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G8gat), .B(G36gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT18), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G64gat), .B(G92gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT26), .B(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313_));
  INV_X1    g112(.A(G183gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT25), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT78), .A3(G183gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT79), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n312_), .A2(KEYINPUT79), .A3(new_n315_), .A4(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n324_), .A2(G169gat), .A3(G176gat), .ZN(new_n325_));
  INV_X1    g124(.A(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT80), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n323_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT23), .B1(new_n314_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT80), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n324_), .B1(G169gat), .B2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(KEYINPUT24), .A4(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n329_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(KEYINPUT82), .A3(new_n333_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n314_), .A2(new_n330_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(new_n332_), .A3(G183gat), .A4(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT22), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G169gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n326_), .A2(KEYINPUT22), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT81), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n350_));
  AOI21_X1  g149(.A(G176gat), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n349_), .A2(new_n351_), .B1(G169gat), .B2(G176gat), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n322_), .A2(new_n339_), .B1(new_n344_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT20), .B1(new_n289_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n323_), .A2(KEYINPUT92), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT24), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n355_), .A2(new_n357_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n340_), .A2(new_n343_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n340_), .A2(KEYINPUT93), .A3(new_n358_), .A4(new_n343_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n355_), .A2(new_n357_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT25), .B(G183gat), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n363_), .A2(new_n364_), .B1(new_n312_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n361_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n334_), .A2(new_n341_), .B1(G169gat), .B2(G176gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n348_), .B(KEYINPUT94), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(G176gat), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n367_), .A2(new_n294_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n354_), .A2(new_n371_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n289_), .B2(new_n353_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n367_), .A2(new_n370_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n285_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n311_), .B1(new_n374_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n322_), .A2(new_n339_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n352_), .A2(new_n344_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n282_), .A2(new_n284_), .A3(KEYINPUT89), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT89), .B1(new_n282_), .B2(new_n284_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT20), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n294_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n373_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n376_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n367_), .A2(new_n294_), .A3(new_n370_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n375_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n310_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n381_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n374_), .A2(new_n380_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT95), .A3(new_n310_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n377_), .A2(new_n379_), .A3(new_n375_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n375_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n311_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(KEYINPUT27), .A3(new_n394_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n306_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n263_), .A2(new_n249_), .A3(new_n261_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(KEYINPUT98), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n245_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n258_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n408_), .B2(KEYINPUT98), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n258_), .A2(new_n413_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n409_), .A2(new_n412_), .B1(new_n266_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n396_), .A2(new_n399_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n265_), .A2(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT99), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT99), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n415_), .A2(new_n416_), .A3(new_n420_), .A4(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT100), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n398_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n373_), .B1(new_n354_), .B2(new_n371_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n425_), .B2(new_n401_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT101), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n426_), .A2(new_n427_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n267_), .A2(new_n265_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n419_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n302_), .A2(new_n305_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n407_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n384_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(new_n242_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G15gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT30), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT31), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n440_), .B(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT102), .B1(new_n435_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT102), .ZN(new_n448_));
  INV_X1    g247(.A(new_n446_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n434_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n418_), .A2(KEYINPUT99), .B1(new_n430_), .B2(new_n431_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n421_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n448_), .B(new_n449_), .C1(new_n452_), .C2(new_n407_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n406_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n431_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n446_), .A3(new_n455_), .A4(new_n434_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G85gat), .B(G92gat), .Z(new_n458_));
  NOR2_X1   g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT7), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n458_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT8), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT10), .B(G99gat), .Z(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(G85gat), .ZN(new_n472_));
  INV_X1    g271(.A(G92gat), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT9), .ZN(new_n474_));
  AOI211_X1 g273(.A(new_n474_), .B(new_n464_), .C1(KEYINPUT9), .C2(new_n458_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n466_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT69), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n471_), .A2(KEYINPUT66), .A3(new_n475_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n466_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n480_), .B(KEYINPUT15), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G232gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n486_), .A2(new_n487_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n482_), .A2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n491_), .A2(new_n488_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G190gat), .B(G218gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT70), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT36), .Z(new_n500_));
  OR2_X1    g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT72), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n495_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n457_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G57gat), .B(G64gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n509_));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n508_), .A2(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n510_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT65), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n477_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n511_), .B(KEYINPUT12), .C1(new_n512_), .C2(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n486_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n515_), .A2(new_n477_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n516_), .B(new_n519_), .C1(new_n520_), .C2(KEYINPUT12), .ZN(new_n521_));
  AND2_X1   g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n516_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n525_), .B2(new_n520_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G176gat), .B(G204gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(KEYINPUT13), .A3(new_n534_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G113gat), .B(G141gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT73), .B(G8gat), .ZN(new_n544_));
  INV_X1    g343(.A(G1gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G1gat), .B(G8gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n548_), .B(KEYINPUT74), .ZN(new_n553_));
  INV_X1    g352(.A(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n487_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n555_), .A3(new_n480_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n556_), .B(new_n480_), .Z(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT76), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n543_), .B1(new_n565_), .B2(KEYINPUT77), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n543_), .A2(KEYINPUT77), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(KEYINPUT76), .B2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XOR2_X1   g372(.A(G183gat), .B(G211gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n556_), .B(new_n576_), .ZN(new_n577_));
  AOI211_X1 g376(.A(new_n571_), .B(new_n575_), .C1(new_n577_), .C2(new_n514_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n514_), .B2(new_n577_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n575_), .B(new_n571_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n515_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n581_), .B2(new_n577_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n540_), .A2(new_n570_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n507_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G1gat), .B1(new_n586_), .B2(new_n455_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n506_), .B(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(new_n584_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT75), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n457_), .A2(new_n569_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n539_), .B(KEYINPUT67), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n545_), .A3(new_n431_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n588_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n598_), .A2(KEYINPUT103), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(KEYINPUT103), .ZN(new_n600_));
  OAI221_X1 g399(.A(new_n587_), .B1(new_n588_), .B2(new_n597_), .C1(new_n599_), .C2(new_n600_), .ZN(G1324gat));
  NAND3_X1  g400(.A1(new_n507_), .A2(new_n406_), .A3(new_n585_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(G8gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n603_), .B1(new_n602_), .B2(G8gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT105), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT39), .ZN(new_n608_));
  INV_X1    g407(.A(new_n606_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT105), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n604_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n611_), .A3(KEYINPUT39), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n596_), .A2(new_n544_), .A3(new_n406_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n608_), .A2(new_n612_), .A3(new_n613_), .A4(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1325gat));
  OAI21_X1  g418(.A(G15gat), .B1(new_n586_), .B2(new_n449_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT41), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n596_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1326gat));
  OAI21_X1  g422(.A(G22gat), .B1(new_n586_), .B2(new_n434_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT42), .ZN(new_n625_));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n596_), .A2(new_n626_), .A3(new_n450_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT107), .Z(G1327gat));
  INV_X1    g428(.A(new_n584_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n540_), .A2(new_n570_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n457_), .A2(new_n632_), .A3(new_n590_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n457_), .B2(new_n590_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT44), .B(new_n631_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G29gat), .B1(new_n639_), .B2(new_n455_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n457_), .A2(new_n569_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n506_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n584_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n540_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n455_), .A2(G29gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n640_), .B1(new_n645_), .B2(new_n646_), .ZN(G1328gat));
  NOR2_X1   g446(.A1(new_n454_), .A2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT109), .B1(new_n645_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT109), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n641_), .A2(new_n651_), .A3(new_n644_), .A4(new_n648_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n650_), .A2(KEYINPUT45), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT45), .B1(new_n650_), .B2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n637_), .A2(new_n406_), .A3(new_n638_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n637_), .A2(KEYINPUT108), .A3(new_n406_), .A4(new_n638_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT110), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT110), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n656_), .A2(new_n657_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(G36gat), .A3(new_n659_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT110), .A3(new_n662_), .A4(new_n655_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1329gat));
  OAI21_X1  g468(.A(G43gat), .B1(new_n639_), .B2(new_n449_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n446_), .A2(new_n437_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n645_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g472(.A(G50gat), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n639_), .A2(new_n674_), .A3(new_n434_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n641_), .A2(new_n450_), .A3(new_n644_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(new_n676_), .ZN(G1331gat));
  NAND4_X1  g476(.A1(new_n507_), .A2(new_n570_), .A3(new_n595_), .A4(new_n630_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n455_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n592_), .A2(new_n539_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n457_), .A2(new_n570_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(KEYINPUT111), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(KEYINPUT111), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n431_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n680_), .B1(new_n687_), .B2(new_n679_), .ZN(G1332gat));
  OAI21_X1  g487(.A(G64gat), .B1(new_n678_), .B2(new_n454_), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n454_), .A2(G64gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n683_), .B2(new_n692_), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n678_), .B2(new_n449_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n449_), .A2(G71gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n683_), .B2(new_n697_), .ZN(G1334gat));
  OAI21_X1  g497(.A(G78gat), .B1(new_n678_), .B2(new_n434_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT50), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n434_), .A2(G78gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n683_), .B2(new_n701_), .ZN(G1335gat));
  NOR2_X1   g501(.A1(new_n633_), .A2(new_n634_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n540_), .A2(new_n570_), .A3(new_n584_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(G85gat), .A3(new_n431_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n457_), .A2(new_n570_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(new_n594_), .A3(new_n643_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n431_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n472_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT114), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT114), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n706_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT115), .Z(G1336gat));
  NAND3_X1  g513(.A1(new_n708_), .A2(new_n473_), .A3(new_n406_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n705_), .A2(new_n406_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n717_), .B2(new_n473_), .ZN(G1337gat));
  AND2_X1   g517(.A1(new_n446_), .A2(new_n467_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n708_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n705_), .A2(new_n446_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT116), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G99gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G99gat), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT117), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n708_), .A2(new_n468_), .A3(new_n450_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n705_), .A2(new_n450_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G106gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT52), .B(new_n468_), .C1(new_n705_), .C2(new_n450_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g532(.A1(new_n590_), .A2(new_n540_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT119), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT118), .B1(new_n569_), .B2(new_n584_), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n569_), .A2(KEYINPUT118), .A3(new_n584_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .A4(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n506_), .B(KEYINPUT37), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(new_n539_), .A3(new_n736_), .A4(new_n737_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT119), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(KEYINPUT54), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(KEYINPUT119), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n563_), .A2(new_n561_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n559_), .B(KEYINPUT121), .Z(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n561_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(new_n543_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n564_), .A2(new_n543_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n751_), .A2(KEYINPUT122), .A3(new_n535_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT122), .B1(new_n751_), .B2(new_n535_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n569_), .A2(new_n534_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n758_), .A2(new_n523_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n523_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n533_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n756_), .B1(new_n761_), .B2(KEYINPUT120), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n761_), .A2(new_n756_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n755_), .B(new_n762_), .C1(KEYINPUT120), .C2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n642_), .B1(new_n754_), .B2(new_n764_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n765_), .A2(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n756_), .ZN(new_n767_));
  AND4_X1   g566(.A1(new_n534_), .A2(new_n767_), .A3(new_n749_), .A4(new_n750_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT58), .B1(new_n768_), .B2(new_n763_), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n769_), .A2(new_n739_), .A3(KEYINPUT123), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT123), .B1(new_n769_), .B2(new_n739_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n768_), .A2(new_n763_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT58), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n765_), .A2(KEYINPUT57), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n766_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n745_), .B1(new_n776_), .B2(new_n584_), .ZN(new_n777_));
  NOR4_X1   g576(.A1(new_n455_), .A2(new_n450_), .A3(new_n449_), .A4(new_n406_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(G113gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n569_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n776_), .A2(new_n584_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n745_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT124), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(KEYINPUT59), .A4(new_n778_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n788_), .B(new_n789_), .C1(new_n777_), .C2(new_n779_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n570_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n782_), .B1(new_n791_), .B2(new_n781_), .ZN(G1340gat));
  INV_X1    g591(.A(G120gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n539_), .B2(KEYINPUT60), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n780_), .B(new_n794_), .C1(KEYINPUT60), .C2(new_n793_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n594_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n793_), .ZN(G1341gat));
  NAND2_X1  g596(.A1(new_n630_), .A2(G127gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n765_), .B(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n630_), .B1(new_n801_), .B2(new_n774_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n630_), .B(new_n778_), .C1(new_n802_), .C2(new_n745_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT125), .ZN(new_n804_));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n799_), .A2(new_n806_), .A3(new_n807_), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n780_), .A2(new_n809_), .A3(new_n642_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n739_), .B1(new_n787_), .B2(new_n790_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n809_), .ZN(G1343gat));
  NOR4_X1   g611(.A1(new_n455_), .A2(new_n406_), .A3(new_n434_), .A4(new_n446_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n785_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n570_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n594_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n212_), .ZN(G1345gat));
  NAND3_X1  g617(.A1(new_n785_), .A2(new_n630_), .A3(new_n813_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  OAI21_X1  g620(.A(G162gat), .B1(new_n814_), .B2(new_n739_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n642_), .A2(new_n221_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n814_), .B2(new_n823_), .ZN(G1347gat));
  NOR3_X1   g623(.A1(new_n450_), .A2(new_n449_), .A3(new_n431_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n406_), .B(new_n825_), .C1(new_n802_), .C2(new_n745_), .ZN(new_n826_));
  OAI21_X1  g625(.A(G169gat), .B1(new_n826_), .B2(new_n570_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n826_), .A2(new_n570_), .A3(new_n369_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT62), .B(G169gat), .C1(new_n826_), .C2(new_n570_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(G1348gat));
  OAI21_X1  g631(.A(G176gat), .B1(new_n826_), .B2(new_n594_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n540_), .A2(new_n327_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n826_), .B2(new_n834_), .ZN(G1349gat));
  NOR3_X1   g634(.A1(new_n826_), .A2(new_n365_), .A3(new_n584_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n777_), .A2(new_n454_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n630_), .A3(new_n825_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n314_), .B2(new_n838_), .ZN(G1350gat));
  OAI21_X1  g638(.A(G190gat), .B1(new_n826_), .B2(new_n739_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n642_), .A2(new_n312_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n826_), .B2(new_n841_), .ZN(G1351gat));
  NOR2_X1   g641(.A1(new_n306_), .A2(new_n446_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(new_n569_), .A3(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT126), .B(G197gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1352gat));
  NAND3_X1  g645(.A1(new_n837_), .A2(new_n595_), .A3(new_n843_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g647(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n785_), .A2(new_n406_), .A3(new_n843_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n584_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT63), .B(G211gat), .Z(new_n852_));
  NAND4_X1  g651(.A1(new_n837_), .A2(new_n630_), .A3(new_n843_), .A4(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1354gat));
  INV_X1    g653(.A(G218gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n850_), .A2(new_n855_), .A3(new_n739_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n843_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n777_), .A2(new_n454_), .A3(new_n506_), .A4(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT127), .ZN(new_n859_));
  AOI21_X1  g658(.A(G218gat), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT127), .B1(new_n850_), .B2(new_n506_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n856_), .B1(new_n860_), .B2(new_n861_), .ZN(G1355gat));
endmodule


