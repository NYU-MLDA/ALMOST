//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n203_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n202_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n210_), .B(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n216_));
  OAI22_X1  g015(.A1(new_n213_), .A2(new_n214_), .B1(new_n216_), .B2(KEYINPUT66), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n202_), .A3(new_n218_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n214_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n212_), .B1(KEYINPUT9), .B2(new_n218_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n206_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n222_), .B(new_n224_), .C1(KEYINPUT9), .C2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n221_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n227_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G230gat), .A2(G233gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT64), .Z(new_n237_));
  NOR2_X1   g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n219_), .A2(new_n221_), .A3(new_n226_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n234_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n234_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n227_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(KEYINPUT12), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT12), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n227_), .A2(new_n244_), .A3(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n238_), .B1(new_n237_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(G204gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G120gat), .B(G148gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT5), .B(G176gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT68), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n246_), .A2(new_n237_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n238_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n253_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT69), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n255_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT98), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G225gat), .A2(G233gat), .ZN(new_n268_));
  AND2_X1   g067(.A1(G127gat), .A2(G134gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G127gat), .A2(G134gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(G113gat), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G127gat), .ZN(new_n272_));
  INV_X1    g071(.A(G134gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G113gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G127gat), .A2(G134gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n271_), .A2(new_n277_), .A3(G120gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(G120gat), .B1(new_n271_), .B2(new_n277_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(KEYINPUT92), .B2(KEYINPUT3), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT92), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n283_), .B(new_n284_), .C1(G141gat), .C2(G148gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT2), .ZN(new_n288_));
  NAND2_X1  g087(.A1(KEYINPUT92), .A2(KEYINPUT3), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n291_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n293_), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n281_), .A2(KEYINPUT89), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n302_), .A2(new_n304_), .B1(G141gat), .B2(G148gat), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n301_), .A2(KEYINPUT91), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT91), .B1(new_n301_), .B2(new_n305_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n280_), .B(new_n294_), .C1(new_n306_), .C2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n305_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n301_), .A2(KEYINPUT91), .A3(new_n305_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n282_), .A2(new_n285_), .B1(KEYINPUT92), .B2(KEYINPUT3), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n291_), .B1(new_n313_), .B2(new_n288_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n311_), .A2(new_n312_), .B1(new_n293_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT86), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n317_));
  INV_X1    g116(.A(G120gat), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n269_), .A2(new_n270_), .A3(G113gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n275_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n271_), .A2(new_n277_), .A3(G120gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(KEYINPUT86), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n268_), .B(new_n308_), .C1(new_n315_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G1gat), .B(G29gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(KEYINPUT4), .B(new_n308_), .C1(new_n315_), .C2(new_n324_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n268_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n278_), .A2(new_n279_), .A3(new_n316_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT86), .B1(new_n321_), .B2(new_n322_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n294_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n338_));
  XOR2_X1   g137(.A(KEYINPUT95), .B(KEYINPUT4), .Z(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT96), .A4(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  AOI211_X1 g143(.A(new_n326_), .B(new_n331_), .C1(new_n334_), .C2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n267_), .B1(new_n345_), .B2(KEYINPUT33), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n334_), .A2(new_n344_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n331_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n325_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT98), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT21), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT93), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(KEYINPUT93), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n356_), .A2(new_n357_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G211gat), .B(G218gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n364_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n365_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n362_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G183gat), .ZN(new_n371_));
  INV_X1    g170(.A(G190gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT23), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(G183gat), .A3(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(G183gat), .B2(G190gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT83), .B(G176gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G169gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT25), .B(G183gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT26), .B(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n375_), .A2(KEYINPUT85), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n373_), .A2(new_n375_), .A3(KEYINPUT85), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT24), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n388_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(KEYINPUT24), .A3(new_n381_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n382_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n370_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n362_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT26), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(G190gat), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n383_), .C1(new_n384_), .C2(new_n398_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n373_), .A2(new_n375_), .B1(new_n389_), .B2(new_n388_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n401_), .A2(KEYINPUT80), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n384_), .A2(new_n398_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n400_), .A4(new_n383_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n402_), .A2(new_n403_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .A4(new_n393_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n379_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT82), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413_));
  INV_X1    g212(.A(G169gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(KEYINPUT22), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n411_), .A2(new_n412_), .A3(new_n415_), .A4(new_n378_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n378_), .B(new_n415_), .C1(new_n413_), .C2(new_n379_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT84), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n386_), .B(new_n387_), .C1(G183gat), .C2(G190gat), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n381_), .A4(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n397_), .B1(new_n409_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n355_), .B1(new_n396_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT18), .B(G64gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G92gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n370_), .B2(new_n395_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n409_), .A2(new_n420_), .A3(new_n397_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n354_), .A3(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n422_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n426_), .B1(new_n422_), .B2(new_n430_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n347_), .A2(KEYINPUT33), .A3(new_n325_), .A4(new_n348_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n344_), .A2(new_n268_), .A3(new_n332_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n308_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT99), .B(new_n308_), .C1(new_n315_), .C2(new_n324_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n333_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n331_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n433_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT100), .B1(new_n352_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n315_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT28), .B1(new_n338_), .B2(KEYINPUT29), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(G22gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n448_), .B(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n370_), .B1(new_n315_), .B2(new_n445_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G50gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G50gat), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n370_), .C1(new_n315_), .C2(new_n445_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n456_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n452_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n451_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n448_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n461_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n459_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n347_), .A2(new_n325_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n331_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n349_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n422_), .A2(new_n430_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n426_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT32), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n354_), .B1(new_n396_), .B2(new_n421_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n428_), .A2(new_n355_), .A3(new_n429_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n470_), .B(new_n474_), .C1(new_n477_), .C2(new_n473_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n433_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n346_), .A4(new_n351_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n443_), .A2(new_n467_), .A3(new_n478_), .A4(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n409_), .A2(new_n420_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n409_), .B2(new_n420_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n409_), .A2(new_n420_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT30), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n490_), .A3(new_n487_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G15gat), .B(G43gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n324_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(new_n496_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n486_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n485_), .A3(new_n500_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n505_), .A3(KEYINPUT88), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n470_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n432_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n422_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT27), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n432_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n467_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n510_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n506_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n467_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT101), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n516_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n512_), .B(KEYINPUT27), .C1(new_n477_), .C2(new_n472_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n467_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT101), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n511_), .A4(new_n506_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n482_), .A2(new_n520_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  INV_X1    g330(.A(G43gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G50gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT70), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n533_), .A2(G50gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(G50gat), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n530_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n534_), .A2(KEYINPUT70), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n533_), .B(new_n457_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n536_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n543_), .A3(KEYINPUT15), .ZN(new_n544_));
  XOR2_X1   g343(.A(KEYINPUT72), .B(G8gat), .Z(new_n545_));
  INV_X1    g344(.A(G1gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT73), .B(G1gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G8gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n540_), .A2(new_n544_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT77), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n552_), .A2(new_n534_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT78), .Z(new_n557_));
  INV_X1    g356(.A(KEYINPUT77), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n540_), .A2(new_n558_), .A3(new_n544_), .A4(new_n552_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n554_), .A2(new_n555_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n552_), .B(new_n534_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(G229gat), .A3(G233gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n414_), .ZN(new_n565_));
  INV_X1    g364(.A(G197gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n560_), .A2(new_n562_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n266_), .A2(new_n529_), .A3(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n540_), .A2(new_n227_), .A3(new_n544_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n239_), .A2(new_n542_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT35), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(KEYINPUT71), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT35), .A3(new_n577_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n581_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G134gat), .ZN(new_n587_));
  INV_X1    g386(.A(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n583_), .A2(new_n584_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT37), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n583_), .A2(new_n594_), .A3(new_n584_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT37), .B1(new_n597_), .B2(new_n590_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n234_), .B(new_n600_), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n552_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT75), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n604_), .B(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n602_), .A2(KEYINPUT17), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT76), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT76), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n617_), .A3(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n599_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n573_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n546_), .A3(new_n470_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT38), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n597_), .A2(new_n590_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n573_), .A2(new_n626_), .A3(new_n615_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n470_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n625_), .B1(new_n630_), .B2(G1gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT103), .B(new_n546_), .C1(new_n629_), .C2(new_n470_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n624_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT104), .B(new_n624_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(new_n518_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n573_), .A2(new_n626_), .A3(new_n638_), .A4(new_n615_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT105), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(KEYINPUT105), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(G8gat), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT106), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n640_), .A2(new_n644_), .A3(G8gat), .A4(new_n641_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(KEYINPUT39), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n622_), .A2(new_n545_), .A3(new_n638_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(KEYINPUT106), .A3(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n646_), .A2(KEYINPUT40), .A3(new_n647_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n629_), .B2(new_n510_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT41), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n622_), .A2(new_n655_), .A3(new_n510_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(new_n467_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n450_), .B1(new_n629_), .B2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT42), .Z(new_n662_));
  NAND3_X1  g461(.A1(new_n622_), .A2(new_n450_), .A3(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n266_), .A2(new_n572_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n482_), .A2(new_n520_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n523_), .A2(new_n528_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n599_), .A3(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n599_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n529_), .B2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n665_), .A2(new_n671_), .A3(new_n675_), .A4(new_n620_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT44), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n511_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n619_), .A2(new_n626_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n573_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n511_), .A2(G29gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT108), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n682_), .B2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n681_), .A2(new_n686_), .A3(new_n638_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT45), .Z(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n677_), .B2(new_n638_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT46), .ZN(G1329gat));
  NAND3_X1  g490(.A1(new_n677_), .A2(G43gat), .A3(new_n506_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT110), .B(G43gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n510_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n682_), .B2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n695_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT47), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n694_), .A2(new_n701_), .A3(new_n695_), .A4(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n681_), .B2(new_n660_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n467_), .A2(new_n457_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n677_), .B2(new_n705_), .ZN(G1331gat));
  NAND2_X1  g505(.A1(new_n264_), .A2(new_n265_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(new_n529_), .A3(new_n571_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n619_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n626_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(G57gat), .A3(new_n470_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT111), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n674_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n470_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1332gat));
  OR3_X1    g515(.A1(new_n713_), .A2(G64gat), .A3(new_n518_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n710_), .A2(new_n638_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G64gat), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT112), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT112), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(KEYINPUT48), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT48), .B1(new_n720_), .B2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(G1333gat));
  NAND2_X1  g523(.A1(new_n710_), .A2(new_n510_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G71gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT49), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n697_), .A2(G71gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n713_), .B2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n710_), .B2(new_n660_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n660_), .A2(new_n730_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT113), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n713_), .B2(new_n734_), .ZN(G1335gat));
  AND2_X1   g534(.A1(new_n708_), .A2(new_n680_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n470_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n707_), .A2(new_n571_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n671_), .A2(new_n675_), .A3(new_n620_), .A4(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n511_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n740_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n736_), .B2(new_n638_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n739_), .A2(new_n518_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n739_), .B2(new_n697_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT114), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n223_), .A3(new_n506_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n746_), .B(new_n747_), .C1(KEYINPUT115), .C2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT115), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(G1338gat));
  AND3_X1   g550(.A1(new_n671_), .A2(new_n675_), .A3(new_n620_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n660_), .A4(new_n738_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n739_), .B2(new_n467_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(G106gat), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n754_), .A2(new_n755_), .A3(new_n758_), .A4(G106gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n736_), .A2(new_n206_), .A3(new_n660_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n757_), .A2(KEYINPUT52), .A3(new_n759_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n762_), .A2(new_n767_), .A3(new_n763_), .A4(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT121), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT57), .ZN(new_n771_));
  INV_X1    g570(.A(new_n626_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n237_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n243_), .A2(new_n773_), .A3(new_n245_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n256_), .A2(KEYINPUT55), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n246_), .A2(new_n777_), .A3(new_n237_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n254_), .A4(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT118), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n775_), .A2(new_n254_), .A3(new_n778_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n258_), .A2(KEYINPUT69), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n247_), .A2(new_n260_), .A3(new_n253_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n781_), .A2(KEYINPUT118), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n780_), .A2(new_n784_), .A3(new_n571_), .A4(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n561_), .A2(new_n557_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n554_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n567_), .B(new_n787_), .C1(new_n788_), .C2(new_n557_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n789_), .A2(new_n570_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n262_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n772_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n771_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n781_), .A2(KEYINPUT118), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n782_), .A2(new_n783_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n571_), .B1(KEYINPUT118), .B2(new_n779_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n791_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n626_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n794_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n785_), .A2(new_n790_), .A3(new_n796_), .A4(new_n779_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n804_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n599_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n802_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n620_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n621_), .A2(new_n707_), .A3(new_n572_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT54), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n621_), .A2(new_n707_), .A3(new_n813_), .A4(new_n572_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT59), .B1(new_n810_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n526_), .A2(new_n470_), .A3(new_n506_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n770_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n809_), .A2(new_n620_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n820_), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n817_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n807_), .B1(new_n794_), .B2(new_n801_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n815_), .B1(new_n823_), .B2(new_n615_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n826_), .B(new_n815_), .C1(new_n823_), .C2(new_n615_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n827_), .A3(new_n818_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n822_), .A2(G113gat), .A3(new_n571_), .A4(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n275_), .B1(new_n828_), .B2(new_n572_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1340gat));
  INV_X1    g631(.A(new_n819_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n816_), .A2(new_n770_), .A3(new_n818_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n829_), .A3(new_n266_), .A4(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G120gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n318_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT122), .B1(new_n318_), .B2(KEYINPUT60), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n828_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n841_), .ZN(G1341gat));
  NAND4_X1  g641(.A1(new_n822_), .A2(G127gat), .A3(new_n615_), .A4(new_n829_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n272_), .B1(new_n828_), .B2(new_n620_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1342gat));
  NAND4_X1  g644(.A1(new_n822_), .A2(G134gat), .A3(new_n599_), .A4(new_n829_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n273_), .B1(new_n828_), .B2(new_n626_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1343gat));
  NOR2_X1   g647(.A1(new_n510_), .A2(new_n467_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n825_), .A2(new_n470_), .A3(new_n827_), .A4(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n638_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n571_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n266_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n619_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  NOR3_X1   g657(.A1(new_n850_), .A2(new_n626_), .A3(new_n638_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT123), .B1(new_n859_), .B2(G162gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n825_), .A2(new_n827_), .A3(new_n849_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n861_), .A2(new_n470_), .A3(new_n772_), .A4(new_n518_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n588_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n674_), .A2(new_n588_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n860_), .A2(new_n864_), .B1(new_n851_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n518_), .A2(new_n470_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n510_), .A2(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n820_), .A2(new_n660_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n571_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n871_), .B2(G169gat), .ZN(new_n872_));
  AOI211_X1 g671(.A(KEYINPUT62), .B(new_n414_), .C1(new_n870_), .C2(new_n571_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n571_), .A2(new_n379_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT124), .ZN(new_n876_));
  OAI22_X1  g675(.A1(new_n872_), .A2(new_n873_), .B1(new_n874_), .B2(new_n876_), .ZN(G1348gat));
  NAND3_X1  g676(.A1(new_n825_), .A2(new_n467_), .A3(new_n827_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n869_), .B1(new_n878_), .B2(KEYINPUT125), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n825_), .A2(new_n880_), .A3(new_n467_), .A4(new_n827_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n879_), .A2(G176gat), .A3(new_n266_), .A4(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n378_), .B1(new_n874_), .B2(new_n707_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1349gat));
  INV_X1    g683(.A(new_n383_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n870_), .A2(new_n885_), .A3(new_n615_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n870_), .A2(KEYINPUT126), .A3(new_n885_), .A4(new_n615_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n879_), .A2(new_n619_), .A3(new_n881_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n371_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n874_), .B2(new_n674_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n870_), .A2(new_n772_), .A3(new_n384_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  NAND4_X1  g694(.A1(new_n825_), .A2(new_n827_), .A3(new_n849_), .A4(new_n868_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n572_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n566_), .ZN(G1352gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n707_), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(G204gat), .Z(G1353gat));
  INV_X1    g699(.A(KEYINPUT127), .ZN(new_n901_));
  NAND2_X1  g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n615_), .A2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n861_), .A2(new_n901_), .A3(new_n868_), .A4(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n903_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT127), .B1(new_n896_), .B2(new_n906_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n904_), .A2(new_n905_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n904_), .B2(new_n907_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1354gat));
  NOR2_X1   g709(.A1(new_n896_), .A2(new_n626_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(G218gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n896_), .A2(new_n674_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(G218gat), .B2(new_n913_), .ZN(G1355gat));
endmodule


