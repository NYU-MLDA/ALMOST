//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  AND3_X1   g003(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT1), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n207_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n210_), .A2(new_n212_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n216_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n218_), .B(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n214_), .B(new_n221_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n219_), .A2(new_n220_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n220_), .B1(new_n219_), .B2(new_n226_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n204_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n219_), .A2(new_n226_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(new_n204_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(KEYINPUT4), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G225gat), .ZN(new_n233_));
  INV_X1    g032(.A(G233gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n236_), .B(new_n204_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT96), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n229_), .A2(new_n231_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n232_), .A2(KEYINPUT96), .A3(new_n235_), .A4(new_n237_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G57gat), .B(G85gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n240_), .A2(new_n242_), .A3(new_n243_), .A4(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n250_), .A2(KEYINPUT99), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT99), .B1(new_n250_), .B2(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n230_), .A2(KEYINPUT86), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n219_), .A2(new_n220_), .A3(new_n226_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT90), .ZN(new_n262_));
  INV_X1    g061(.A(G204gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(G197gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(G197gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(KEYINPUT89), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT89), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n269_), .B2(G197gat), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n261_), .B(new_n264_), .C1(new_n270_), .C2(new_n262_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n269_), .A2(G197gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT88), .ZN(new_n273_));
  INV_X1    g072(.A(G197gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(G204gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n263_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT21), .B1(new_n272_), .B2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G211gat), .B(G218gat), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n264_), .B1(new_n270_), .B2(new_n262_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT21), .A3(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT87), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(G228gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(G228gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n234_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n281_), .A2(new_n283_), .B1(new_n230_), .B2(KEYINPUT29), .ZN(new_n292_));
  OAI22_X1  g091(.A1(new_n260_), .A2(new_n291_), .B1(new_n292_), .B2(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G78gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n289_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n227_), .A2(new_n228_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n257_), .ZN(new_n297_));
  INV_X1    g096(.A(G78gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n230_), .A2(KEYINPUT29), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n284_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n289_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n294_), .A2(G106gat), .A3(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(G106gat), .B1(new_n294_), .B2(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n256_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n296_), .A2(new_n257_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT28), .B(G22gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G50gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n306_), .B(new_n308_), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G106gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n293_), .A2(G78gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n298_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n294_), .A2(new_n302_), .A3(G106gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT91), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n305_), .A2(new_n310_), .A3(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n256_), .B(new_n309_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT80), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT78), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n325_), .B2(KEYINPUT23), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n327_));
  AOI211_X1 g126(.A(KEYINPUT80), .B(new_n327_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n321_), .A2(KEYINPUT23), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT81), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(KEYINPUT23), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT80), .ZN(new_n334_));
  INV_X1    g133(.A(new_n329_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n325_), .A2(new_n320_), .A3(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  INV_X1    g137(.A(new_n331_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT79), .Z(new_n345_));
  NAND3_X1  g144(.A1(new_n332_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(new_n341_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT25), .B(G183gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT26), .B(G190gat), .ZN(new_n351_));
  AOI211_X1 g150(.A(new_n347_), .B(new_n349_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n325_), .A2(new_n327_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n346_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT30), .ZN(new_n357_));
  XOR2_X1   g156(.A(G15gat), .B(G43gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n346_), .A2(new_n366_), .A3(new_n355_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n363_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n357_), .A2(new_n365_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n357_), .A2(new_n367_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT83), .B(new_n369_), .C1(new_n370_), .C2(new_n365_), .ZN(new_n371_));
  XOR2_X1   g170(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n204_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n371_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n319_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n371_), .B(new_n373_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n255_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT100), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n356_), .B2(new_n284_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n284_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n353_), .A2(new_n354_), .A3(new_n339_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n344_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n337_), .A2(new_n352_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n383_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n337_), .A2(KEYINPUT93), .A3(new_n352_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT93), .B1(new_n337_), .B2(new_n352_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n388_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n284_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n346_), .A2(new_n355_), .A3(new_n386_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT20), .ZN(new_n397_));
  INV_X1    g196(.A(new_n383_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n391_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n380_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n380_), .B(new_n406_), .C1(new_n391_), .C2(new_n399_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT27), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n397_), .A2(new_n398_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n356_), .A2(new_n284_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n386_), .B(new_n388_), .C1(new_n393_), .C2(new_n392_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(KEYINPUT20), .A3(new_n383_), .A4(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n413_), .A3(new_n405_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n407_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n406_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT95), .A3(new_n414_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT95), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n410_), .A2(new_n413_), .A3(new_n421_), .A4(new_n405_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT101), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT101), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n419_), .A2(new_n425_), .A3(new_n420_), .A4(new_n422_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n416_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n317_), .A2(new_n318_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n419_), .A2(new_n422_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n252_), .B(KEYINPUT33), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n251_), .B1(new_n241_), .B2(new_n235_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n232_), .A2(new_n237_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n235_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n400_), .A2(KEYINPUT32), .A3(new_n405_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n250_), .A2(new_n252_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT98), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n435_), .B(new_n436_), .C1(new_n417_), .C2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n428_), .B1(new_n434_), .B2(new_n439_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n379_), .A2(new_n427_), .B1(new_n440_), .B2(new_n377_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT73), .B(G22gat), .ZN(new_n442_));
  INV_X1    g241(.A(G15gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G1gat), .ZN(new_n445_));
  INV_X1    g244(.A(G8gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT14), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G8gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n448_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G57gat), .ZN(new_n452_));
  INV_X1    g251(.A(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G57gat), .A2(G64gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT66), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT66), .B1(new_n454_), .B2(new_n455_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT11), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G71gat), .B(G78gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n456_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n461_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n464_), .B2(new_n456_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n460_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n451_), .B(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(G231gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G127gat), .B(G155gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G211gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT16), .B(G183gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT74), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT17), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(KEYINPUT17), .B2(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n473_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT69), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G85gat), .B(G92gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT10), .B(G99gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n311_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(G85gat), .A3(G92gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n489_), .A2(new_n491_), .A3(new_n497_), .ZN(new_n498_));
  OR3_X1    g297(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n499_), .A2(new_n494_), .A3(new_n496_), .A4(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G85gat), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n505_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n501_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT8), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n487_), .A2(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n507_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n501_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n498_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G29gat), .B(G36gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(G29gat), .B(G36gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT15), .B1(new_n519_), .B2(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n486_), .B1(new_n516_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n498_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n513_), .A2(new_n514_), .A3(new_n501_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n514_), .B1(new_n513_), .B2(new_n501_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n523_), .B(new_n524_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT69), .ZN(new_n534_));
  INV_X1    g333(.A(new_n523_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n516_), .A2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n528_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT35), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n528_), .A2(new_n534_), .A3(new_n544_), .A4(new_n536_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(new_n538_), .A3(KEYINPUT35), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT70), .B1(new_n542_), .B2(new_n543_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n541_), .A2(KEYINPUT36), .A3(new_n548_), .A4(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n541_), .A2(new_n548_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(KEYINPUT71), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557_));
  INV_X1    g356(.A(new_n554_), .ZN(new_n558_));
  AOI211_X1 g357(.A(new_n557_), .B(new_n558_), .C1(new_n541_), .C2(new_n548_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n553_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n553_), .B(new_n561_), .C1(new_n556_), .C2(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n441_), .A2(new_n485_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n451_), .A2(new_n535_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n448_), .B(new_n449_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n533_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT75), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n569_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT76), .ZN(new_n573_));
  INV_X1    g372(.A(new_n570_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n567_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n451_), .A2(new_n535_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n567_), .A2(new_n569_), .A3(new_n578_), .A4(new_n571_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  INV_X1    g380(.A(G141gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT77), .B(G113gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n573_), .A2(new_n577_), .A3(new_n579_), .A4(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT67), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  OAI22_X1  g390(.A1(new_n516_), .A2(new_n470_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n516_), .A2(new_n470_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT64), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n591_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n467_), .A2(new_n469_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n590_), .A2(new_n591_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n532_), .A3(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .A4(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n596_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n593_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n516_), .A2(new_n470_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(G204gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT5), .B(G176gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n601_), .A2(new_n605_), .A3(new_n612_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n611_), .A2(KEYINPUT13), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT13), .B1(new_n611_), .B2(new_n613_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT68), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n566_), .A2(new_n589_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n445_), .A3(new_n255_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n376_), .A2(new_n378_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n424_), .A2(new_n426_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n255_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n416_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .A4(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n434_), .A2(new_n439_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n377_), .A3(new_n319_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n560_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n553_), .B(KEYINPUT102), .C1(new_n556_), .C2(new_n559_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n485_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n616_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n589_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n629_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n445_), .B1(new_n644_), .B2(new_n255_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT104), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT104), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n621_), .B1(new_n646_), .B2(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(new_n427_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n619_), .A2(new_n446_), .A3(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n629_), .A2(new_n635_), .A3(new_n638_), .A4(new_n649_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G8gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT105), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n655_), .A3(G8gat), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n653_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n654_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n650_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1325gat));
  NAND3_X1  g460(.A1(new_n619_), .A2(new_n443_), .A3(new_n375_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n643_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n375_), .B1(new_n663_), .B2(new_n641_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G15gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT106), .B(KEYINPUT107), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(G15gat), .A3(new_n666_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(KEYINPUT41), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n668_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n662_), .B1(new_n670_), .B2(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n428_), .B(KEYINPUT108), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n619_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n677_), .A2(new_n673_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT42), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(KEYINPUT42), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NOR3_X1   g480(.A1(new_n441_), .A2(new_n637_), .A3(new_n636_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n633_), .A2(new_n484_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT110), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n255_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n565_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT109), .B(new_n692_), .C1(new_n441_), .C2(new_n688_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n636_), .A2(new_n484_), .A3(new_n637_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n691_), .A2(KEYINPUT44), .A3(new_n693_), .A4(new_n694_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(G29gat), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n687_), .B1(new_n699_), .B2(new_n255_), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n698_), .A2(new_n649_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n697_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n682_), .A2(new_n705_), .A3(new_n649_), .A4(new_n684_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT45), .Z(new_n709_));
  OAI211_X1 g508(.A(new_n703_), .B(new_n704_), .C1(new_n707_), .C2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n697_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n698_), .A2(new_n649_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G36gat), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(new_n701_), .A3(new_n702_), .A4(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n710_), .A2(new_n715_), .ZN(G1329gat));
  NAND3_X1  g515(.A1(new_n698_), .A2(G43gat), .A3(new_n375_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n685_), .A2(new_n377_), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n711_), .A2(new_n717_), .B1(G43gat), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n697_), .A2(new_n428_), .A3(new_n698_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G50gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n674_), .A2(G50gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT112), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n685_), .B2(new_n724_), .ZN(G1331gat));
  NOR3_X1   g524(.A1(new_n441_), .A2(new_n618_), .A3(new_n589_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n635_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(new_n452_), .A3(new_n624_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n616_), .A2(new_n589_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n566_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n255_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n452_), .B2(new_n732_), .ZN(G1332gat));
  NAND3_X1  g532(.A1(new_n731_), .A2(new_n453_), .A3(new_n649_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G64gat), .B1(new_n727_), .B2(new_n427_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT48), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT48), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(G1333gat));
  OR3_X1    g537(.A1(new_n730_), .A2(G71gat), .A3(new_n377_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n726_), .A2(new_n635_), .A3(new_n375_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(G71gat), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G71gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n727_), .B2(new_n674_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(KEYINPUT114), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(KEYINPUT114), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n674_), .A2(G78gat), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT115), .ZN(new_n752_));
  OAI22_X1  g551(.A1(new_n749_), .A2(new_n750_), .B1(new_n730_), .B2(new_n752_), .ZN(G1335gat));
  AND2_X1   g552(.A1(new_n726_), .A2(new_n684_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754_), .B2(new_n255_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n691_), .A2(new_n693_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n729_), .A2(new_n485_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT116), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n624_), .A2(new_n502_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n760_), .B2(new_n761_), .ZN(G1336gat));
  AOI21_X1  g561(.A(G92gat), .B1(new_n754_), .B2(new_n649_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n427_), .A2(new_n503_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n760_), .B2(new_n764_), .ZN(G1337gat));
  NOR2_X1   g564(.A1(new_n377_), .A2(new_n490_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n754_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n759_), .A2(new_n377_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n493_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n767_), .C1(new_n768_), .C2(new_n493_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n754_), .A2(new_n311_), .A3(new_n428_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n691_), .A2(new_n428_), .A3(new_n693_), .A4(new_n758_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G106gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n649_), .A2(new_n624_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n376_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n592_), .A2(new_n600_), .A3(new_n593_), .A4(new_n597_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n602_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n612_), .B1(new_n788_), .B2(new_n601_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n592_), .A2(new_n600_), .A3(new_n593_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(new_n786_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(KEYINPUT56), .A4(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n589_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n602_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT55), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n787_), .A2(new_n602_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n610_), .B(new_n792_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n792_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(KEYINPUT117), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n794_), .A2(new_n802_), .A3(new_n613_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n611_), .A2(new_n613_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n571_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n567_), .A2(new_n569_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n805_), .B(new_n585_), .C1(new_n806_), .C2(new_n571_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n588_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n803_), .A2(new_n809_), .B1(new_n632_), .B2(new_n631_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n785_), .B1(new_n810_), .B2(KEYINPUT57), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n785_), .A3(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n803_), .A2(new_n809_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n633_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(KEYINPUT118), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n818_), .B1(new_n810_), .B2(KEYINPUT57), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n812_), .A2(new_n813_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n800_), .A2(new_n801_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n613_), .A3(new_n808_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n821_), .A2(new_n613_), .A3(new_n826_), .A4(new_n808_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n565_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n484_), .B1(new_n820_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n565_), .A2(new_n485_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n637_), .A3(new_n616_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT54), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n830_), .A2(new_n833_), .A3(new_n637_), .A4(new_n616_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n784_), .B1(new_n829_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n589_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n828_), .B(KEYINPUT121), .C1(new_n810_), .C2(KEYINPUT57), .ZN(new_n840_));
  AND4_X1   g639(.A1(new_n785_), .A2(new_n814_), .A3(new_n633_), .A4(KEYINPUT57), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n811_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n815_), .A2(new_n816_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT121), .B1(new_n843_), .B2(new_n828_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n485_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT122), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n847_), .B(new_n485_), .C1(new_n842_), .C2(new_n844_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n835_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n784_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n589_), .A2(G113gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n839_), .B1(new_n853_), .B2(new_n854_), .ZN(G1340gat));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n617_), .A3(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT60), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n616_), .B2(G120gat), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n838_), .B(new_n859_), .C1(new_n858_), .C2(G120gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1341gat));
  AND4_X1   g660(.A1(G127gat), .A2(new_n851_), .A3(new_n484_), .A4(new_n852_), .ZN(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n837_), .B2(new_n485_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT123), .B(new_n863_), .C1(new_n837_), .C2(new_n485_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n862_), .A2(new_n868_), .ZN(G1342gat));
  AOI21_X1  g668(.A(G134gat), .B1(new_n838_), .B2(new_n634_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n565_), .A2(G134gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n853_), .B2(new_n871_), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n817_), .A2(new_n819_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n873_), .B(new_n828_), .C1(new_n811_), .C2(new_n841_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n836_), .B1(new_n874_), .B2(new_n485_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n378_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n781_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n637_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n582_), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n876_), .A2(new_n617_), .A3(new_n781_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g680(.A1(new_n877_), .A2(new_n485_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n877_), .A2(new_n885_), .A3(new_n688_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n876_), .A2(new_n634_), .A3(new_n781_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(G162gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT124), .B(new_n885_), .C1(new_n877_), .C2(new_n633_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n889_), .B2(new_n890_), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n427_), .A2(new_n255_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n375_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n675_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n849_), .A2(new_n589_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n895_), .A2(G169gat), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(G169gat), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n849_), .A2(new_n589_), .A3(new_n342_), .A4(new_n894_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n900_), .A2(new_n896_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n899_), .B2(new_n901_), .ZN(G1348gat));
  AND2_X1   g701(.A1(new_n849_), .A2(new_n894_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G176gat), .B1(new_n903_), .B2(new_n636_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n875_), .A2(new_n428_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n893_), .A2(new_n618_), .A3(new_n343_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1349gat));
  NOR2_X1   g706(.A1(new_n485_), .A2(new_n350_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n905_), .A2(new_n484_), .A3(new_n375_), .A4(new_n892_), .ZN(new_n909_));
  INV_X1    g708(.A(G183gat), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n903_), .A2(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1350gat));
  NAND2_X1  g710(.A1(new_n903_), .A2(new_n565_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G190gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n903_), .A2(new_n634_), .A3(new_n351_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1351gat));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  INV_X1    g715(.A(new_n378_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(new_n892_), .C1(new_n829_), .C2(new_n836_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n637_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n916_), .B1(new_n919_), .B2(G197gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(G197gat), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT126), .B(new_n274_), .C1(new_n918_), .C2(new_n637_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(G1352gat));
  NOR2_X1   g722(.A1(new_n918_), .A2(new_n618_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n269_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n924_), .B2(new_n263_), .ZN(G1353gat));
  OAI22_X1  g725(.A1(new_n918_), .A2(new_n485_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT63), .B(G211gat), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n876_), .A2(new_n484_), .A3(new_n892_), .A4(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n927_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n927_), .B2(new_n929_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1354gat));
  INV_X1    g732(.A(G218gat), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n918_), .A2(new_n934_), .A3(new_n688_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n876_), .A2(new_n634_), .A3(new_n892_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n934_), .ZN(G1355gat));
endmodule


