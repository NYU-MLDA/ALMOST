//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_;
  INV_X1    g000(.A(KEYINPUT26), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(G183gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT25), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT26), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT103), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT103), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT23), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n222_), .A2(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT104), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n211_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n231_), .A3(new_n212_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n214_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n222_), .A2(new_n224_), .B1(new_n204_), .B2(new_n208_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n228_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n214_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G169gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(new_n237_), .B2(new_n212_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n222_), .A2(new_n224_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n204_), .A2(new_n208_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n241_), .A3(KEYINPUT104), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n220_), .A2(new_n227_), .B1(new_n235_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT98), .ZN(new_n244_));
  INV_X1    g043(.A(G211gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G218gat), .ZN(new_n246_));
  INV_X1    g045(.A(G218gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(G211gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(G211gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(G218gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT98), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT21), .ZN(new_n253_));
  INV_X1    g052(.A(G204gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G197gat), .ZN(new_n255_));
  INV_X1    g054(.A(G197gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G204gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n253_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n252_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT99), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n249_), .A2(KEYINPUT99), .A3(new_n258_), .A4(new_n252_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n255_), .A2(new_n257_), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n264_));
  AOI22_X1  g063(.A1(new_n249_), .A2(new_n252_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n257_), .A2(KEYINPUT96), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n255_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n257_), .A2(KEYINPUT96), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT21), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n261_), .A2(new_n262_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT20), .B1(new_n243_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT81), .B1(new_n208_), .B2(KEYINPUT26), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n202_), .A3(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n208_), .A2(KEYINPUT80), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G190gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT26), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT25), .B(G183gat), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n275_), .A2(new_n279_), .A3(KEYINPUT82), .A4(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n225_), .B1(G169gat), .B2(G176gat), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT83), .B1(new_n286_), .B2(new_n213_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n214_), .A2(KEYINPUT24), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n226_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n227_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n230_), .A2(KEYINPUT84), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT22), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n211_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n298_));
  AOI21_X1  g097(.A(G176gat), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n229_), .A2(new_n298_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n294_), .A2(new_n296_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(new_n211_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n276_), .A2(new_n278_), .A3(new_n204_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n239_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n214_), .A3(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n270_), .A2(new_n293_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT19), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n271_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n261_), .A2(new_n262_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n265_), .A2(new_n269_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n291_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n214_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n302_), .B2(new_n299_), .ZN(new_n316_));
  OAI22_X1  g115(.A1(new_n311_), .A2(new_n313_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n210_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n218_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n227_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n234_), .B2(new_n233_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n261_), .A2(new_n262_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n312_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT20), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n309_), .B1(new_n318_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n310_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n309_), .B1(new_n271_), .B2(new_n307_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n235_), .A2(new_n242_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n323_), .A2(new_n321_), .A3(new_n312_), .A4(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT105), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n309_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n270_), .A2(KEYINPUT105), .A3(new_n321_), .A4(new_n335_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .A4(new_n317_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n334_), .A2(new_n331_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n334_), .A2(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n332_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n334_), .A2(new_n342_), .A3(new_n331_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n333_), .A2(new_n345_), .B1(new_n349_), .B2(new_n344_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT86), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT87), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n353_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n355_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n293_), .A2(KEYINPUT30), .A3(new_n306_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n364_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  INV_X1    g168(.A(G134gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G127gat), .ZN(new_n371_));
  INV_X1    g170(.A(G127gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G134gat), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT89), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT89), .B1(new_n371_), .B2(new_n373_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT89), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n372_), .A2(G134gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n370_), .A2(G127gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n369_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT89), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n376_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT31), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT90), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n366_), .A2(new_n368_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT91), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT90), .B1(new_n385_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT91), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n366_), .A2(new_n391_), .A3(new_n368_), .A4(new_n386_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n350_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT94), .A3(KEYINPUT1), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT94), .B1(new_n402_), .B2(KEYINPUT1), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT93), .ZN(new_n407_));
  INV_X1    g206(.A(G155gat), .ZN(new_n408_));
  INV_X1    g207(.A(G162gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT93), .B1(G155gat), .B2(G162gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(G155gat), .A3(G162gat), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n401_), .B1(new_n406_), .B2(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n399_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT2), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n397_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n416_), .A2(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n374_), .A2(new_n375_), .A3(new_n369_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n381_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n426_));
  OAI22_X1  g225(.A1(new_n415_), .A2(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n402_), .A2(KEYINPUT1), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n403_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n400_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n423_), .A2(new_n410_), .A3(new_n411_), .A4(new_n402_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n383_), .A4(new_n376_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n427_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n427_), .A2(KEYINPUT4), .A3(new_n435_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT106), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n427_), .A2(new_n435_), .A3(KEYINPUT106), .A4(KEYINPUT4), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n434_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n384_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n436_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT107), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT107), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n450_), .B(new_n447_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n437_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G1gat), .B(G29gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT0), .ZN(new_n454_));
  INV_X1    g253(.A(G57gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G85gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n437_), .B(new_n457_), .C1(new_n449_), .C2(new_n451_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OR3_X1    g260(.A1(new_n443_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT28), .B1(new_n443_), .B2(KEYINPUT29), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G22gat), .B(G50gat), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G228gat), .ZN(new_n468_));
  INV_X1    g267(.A(G233gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n443_), .A2(KEYINPUT29), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n324_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n443_), .A2(KEYINPUT95), .A3(KEYINPUT29), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n324_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT95), .B1(new_n443_), .B2(KEYINPUT29), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT100), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n470_), .B1(new_n323_), .B2(new_n312_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .A4(new_n474_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n473_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT101), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n467_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  AOI211_X1 g286(.A(new_n487_), .B(new_n473_), .C1(new_n477_), .C2(new_n482_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT102), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n473_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n491_));
  AOI211_X1 g290(.A(new_n478_), .B(new_n491_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n492_), .A2(new_n270_), .A3(new_n470_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n481_), .B1(new_n493_), .B2(new_n479_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n482_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n490_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n487_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT102), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n483_), .A2(new_n485_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .A4(new_n467_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n467_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n483_), .A2(new_n484_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n489_), .A2(new_n500_), .A3(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n396_), .A2(new_n461_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n459_), .A2(new_n460_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n508_), .A3(new_n350_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT110), .ZN(new_n510_));
  INV_X1    g309(.A(new_n506_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n331_), .B1(new_n334_), .B2(new_n342_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n343_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n427_), .A2(new_n435_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT108), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n457_), .B1(new_n515_), .B2(new_n446_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n445_), .A2(new_n436_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n442_), .A2(KEYINPUT109), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT109), .B1(new_n442_), .B2(new_n517_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n513_), .B(new_n520_), .C1(new_n460_), .C2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n460_), .A2(new_n521_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n327_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n334_), .A2(new_n342_), .A3(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n511_), .B1(new_n524_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT110), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n506_), .A2(new_n508_), .A3(new_n350_), .A4(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n510_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n534_));
  OR3_X1    g333(.A1(new_n394_), .A2(KEYINPUT92), .A3(new_n395_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT92), .B1(new_n394_), .B2(new_n395_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n507_), .B1(new_n534_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G169gat), .B(G197gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544_));
  INV_X1    g343(.A(G1gat), .ZN(new_n545_));
  INV_X1    g344(.A(G8gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G8gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G29gat), .B(G36gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT78), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n550_), .A2(new_n553_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT78), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n558_), .B2(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n553_), .B(KEYINPUT15), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n550_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n561_), .B1(new_n564_), .B2(new_n556_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n543_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT79), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT79), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n568_), .B(new_n543_), .C1(new_n562_), .C2(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n562_), .A2(new_n565_), .A3(new_n543_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n539_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT68), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G85gat), .B(G92gat), .Z(new_n581_));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT6), .Z(new_n583_));
  OR3_X1    g382(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n581_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT8), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT65), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(G85gat), .B2(G92gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT64), .B(G92gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(new_n593_), .B2(G85gat), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT66), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n597_));
  INV_X1    g396(.A(G106gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT10), .B(G99gat), .Z(new_n599_));
  AOI21_X1  g398(.A(new_n583_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n588_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n604_));
  XOR2_X1   g403(.A(G71gat), .B(G78gat), .Z(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n604_), .A2(new_n605_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT67), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT67), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n602_), .A2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(G230gat), .A3(G233gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n610_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n614_), .A2(KEYINPUT12), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n614_), .A2(KEYINPUT12), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n617_), .B(new_n618_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n580_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n611_), .A2(new_n612_), .B1(new_n609_), .B2(new_n602_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n621_), .B(new_n580_), .C1(new_n623_), .C2(new_n617_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT13), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n623_), .A2(new_n617_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n621_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n579_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G190gat), .B(G218gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT71), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT72), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT36), .Z(new_n639_));
  AND2_X1   g438(.A1(new_n602_), .A2(new_n563_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT34), .Z(new_n642_));
  INV_X1    g441(.A(KEYINPUT35), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT70), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n602_), .B2(new_n553_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT69), .B(new_n645_), .C1(new_n602_), .C2(new_n553_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n642_), .A2(new_n643_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n648_), .B(new_n649_), .C1(new_n640_), .C2(new_n646_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT73), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n639_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT73), .B1(new_n651_), .B2(new_n652_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n638_), .A2(KEYINPUT36), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n651_), .A2(new_n658_), .A3(new_n652_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(G231gat), .A2(G233gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n550_), .B(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(new_n609_), .ZN(new_n663_));
  XOR2_X1   g462(.A(G127gat), .B(G155gat), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT16), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G183gat), .B(G211gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT17), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n663_), .A2(KEYINPUT76), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT76), .B1(new_n663_), .B2(new_n669_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n667_), .A2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n663_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n660_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n633_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n574_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G1gat), .B1(new_n678_), .B2(new_n508_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n506_), .A2(new_n508_), .A3(new_n350_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n529_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n461_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n447_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT107), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n685_), .A2(KEYINPUT33), .A3(new_n437_), .A4(new_n457_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n460_), .A2(new_n521_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n513_), .A4(new_n520_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n683_), .A2(new_n688_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n681_), .A2(new_n532_), .B1(new_n689_), .B2(new_n511_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n537_), .B1(new_n690_), .B2(new_n510_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n680_), .B(new_n572_), .C1(new_n691_), .C2(new_n507_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT111), .B1(new_n539_), .B2(new_n573_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n633_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n695_));
  OAI211_X1 g494(.A(new_n659_), .B(new_n695_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT75), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n653_), .A2(new_n639_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n659_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT37), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n699_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n674_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT77), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n694_), .A2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n461_), .B(KEYINPUT112), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n545_), .A3(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT38), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT38), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n679_), .B1(new_n710_), .B2(new_n711_), .ZN(G1324gat));
  INV_X1    g511(.A(new_n350_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n546_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n678_), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT39), .B(new_n546_), .C1(new_n715_), .C2(new_n713_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT39), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n713_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G8gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT40), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n714_), .B(KEYINPUT40), .C1(new_n719_), .C2(new_n716_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1325gat));
  OAI21_X1  g523(.A(G15gat), .B1(new_n678_), .B2(new_n538_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT41), .Z(new_n726_));
  INV_X1    g525(.A(G15gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n707_), .A2(new_n727_), .A3(new_n537_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1326gat));
  INV_X1    g528(.A(G22gat), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n506_), .B(KEYINPUT113), .Z(new_n731_));
  NAND3_X1  g530(.A1(new_n707_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n715_), .A2(new_n731_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G22gat), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(KEYINPUT42), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(KEYINPUT42), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1327gat));
  NOR2_X1   g536(.A1(KEYINPUT114), .A2(KEYINPUT44), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(new_n704_), .C1(new_n691_), .C2(new_n507_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n699_), .A2(new_n703_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n539_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n632_), .A2(new_n572_), .A3(new_n674_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n739_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n745_), .B(new_n738_), .C1(new_n741_), .C2(new_n743_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n708_), .ZN(new_n750_));
  INV_X1    g549(.A(G29gat), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n660_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n674_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n694_), .A2(new_n461_), .A3(new_n755_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n749_), .A2(new_n752_), .B1(new_n751_), .B2(new_n756_), .ZN(G1328gat));
  XOR2_X1   g556(.A(KEYINPUT115), .B(KEYINPUT46), .Z(new_n758_));
  INV_X1    g557(.A(G36gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n749_), .B2(new_n713_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n692_), .A2(new_n693_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n350_), .A2(G36gat), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n632_), .A3(new_n755_), .A4(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n758_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n763_), .B(KEYINPUT45), .ZN(new_n767_));
  INV_X1    g566(.A(new_n758_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n747_), .A2(new_n748_), .A3(new_n350_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n767_), .B(new_n768_), .C1(new_n769_), .C2(new_n759_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(new_n770_), .ZN(G1329gat));
  XOR2_X1   g570(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(G43gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n694_), .A2(new_n537_), .A3(new_n755_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n395_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n776_), .B2(new_n393_), .ZN(new_n777_));
  AOI221_X4 g576(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .C1(new_n749_), .C2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n749_), .A2(new_n777_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n774_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n772_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n778_), .A2(new_n781_), .ZN(G1330gat));
  INV_X1    g581(.A(G50gat), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n511_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n694_), .A2(new_n731_), .A3(new_n755_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n749_), .A2(new_n784_), .B1(new_n783_), .B2(new_n785_), .ZN(G1331gat));
  NOR2_X1   g585(.A1(new_n632_), .A2(new_n572_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n691_), .B2(new_n507_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n706_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n455_), .A3(new_n708_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n788_), .A2(new_n508_), .A3(new_n676_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n455_), .B2(new_n792_), .ZN(G1332gat));
  INV_X1    g592(.A(G64gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n794_), .A3(new_n713_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n788_), .A2(new_n676_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n713_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(G64gat), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT48), .B(new_n794_), .C1(new_n797_), .C2(new_n713_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT117), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n795_), .B(new_n803_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1333gat));
  INV_X1    g604(.A(G71gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n797_), .B2(new_n537_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT49), .Z(new_n808_));
  NAND3_X1  g607(.A1(new_n790_), .A2(new_n806_), .A3(new_n537_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1334gat));
  INV_X1    g609(.A(G78gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n797_), .B2(new_n731_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT50), .Z(new_n813_));
  NAND3_X1  g612(.A1(new_n790_), .A2(new_n811_), .A3(new_n731_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1335gat));
  NAND2_X1  g614(.A1(new_n787_), .A2(new_n674_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818_), .B2(new_n508_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n788_), .A2(new_n754_), .ZN(new_n820_));
  INV_X1    g619(.A(G85gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n708_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(G1336gat));
  AOI21_X1  g622(.A(G92gat), .B1(new_n820_), .B2(new_n713_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n713_), .A2(new_n593_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(KEYINPUT118), .Z(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n817_), .B2(new_n826_), .ZN(G1337gat));
  OAI211_X1 g626(.A(new_n820_), .B(new_n599_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n818_), .A2(new_n538_), .ZN(new_n829_));
  INV_X1    g628(.A(G99gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n598_), .A3(new_n506_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n817_), .A2(new_n506_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G106gat), .ZN(new_n836_));
  AOI211_X1 g635(.A(KEYINPUT52), .B(new_n598_), .C1(new_n817_), .C2(new_n506_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT53), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n840_), .B(new_n833_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1339gat));
  NAND2_X1  g641(.A1(new_n572_), .A2(new_n624_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n618_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(G230gat), .A3(G233gat), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n621_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n614_), .B(KEYINPUT12), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n848_), .A2(KEYINPUT55), .A3(new_n617_), .A4(new_n618_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n579_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(KEYINPUT56), .A3(new_n579_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n843_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n629_), .A2(new_n624_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n564_), .A2(new_n556_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT119), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n561_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n559_), .A2(new_n561_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n543_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n567_), .A2(new_n569_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n856_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n660_), .B1(new_n855_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n862_), .A2(new_n624_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n854_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT56), .B1(new_n850_), .B2(new_n579_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n867_), .B(KEYINPUT58), .C1(new_n868_), .C2(new_n869_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n704_), .A3(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT57), .B(new_n660_), .C1(new_n855_), .C2(new_n863_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n866_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n674_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n572_), .B1(new_n626_), .B2(new_n631_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n878_), .B(new_n675_), .C1(new_n699_), .C2(new_n703_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT54), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n750_), .A2(new_n506_), .A3(new_n396_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(G113gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n572_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT59), .B1(new_n881_), .B2(KEYINPUT120), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n883_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n881_), .B(new_n882_), .C1(KEYINPUT120), .C2(KEYINPUT59), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n573_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n886_), .B1(new_n890_), .B2(new_n885_), .ZN(G1340gat));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n892_));
  INV_X1    g691(.A(G120gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n633_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n884_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n632_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n893_), .ZN(G1341gat));
  NAND3_X1  g697(.A1(new_n884_), .A2(new_n372_), .A3(new_n675_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n674_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n372_), .ZN(G1342gat));
  AOI21_X1  g700(.A(G134gat), .B1(new_n884_), .B2(new_n753_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n888_), .A2(new_n889_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT121), .B(G134gat), .Z(new_n904_));
  NOR2_X1   g703(.A1(new_n742_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n903_), .B2(new_n905_), .ZN(G1343gat));
  NOR4_X1   g705(.A1(new_n750_), .A2(new_n537_), .A3(new_n511_), .A4(new_n713_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n881_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n573_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n632_), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(G148gat), .Z(G1345gat));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n908_), .B2(new_n674_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n881_), .A2(KEYINPUT122), .A3(new_n675_), .A4(new_n907_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n908_), .B2(new_n742_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n753_), .A2(new_n409_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n908_), .B2(new_n921_), .ZN(G1347gat));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n750_), .A2(new_n537_), .A3(new_n713_), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT123), .Z(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n731_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n881_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n573_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n923_), .B1(new_n928_), .B2(new_n211_), .ZN(new_n929_));
  OAI211_X1 g728(.A(KEYINPUT62), .B(G169gat), .C1(new_n927_), .C2(new_n573_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n237_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(G1348gat));
  INV_X1    g731(.A(new_n927_), .ZN(new_n933_));
  AOI21_X1  g732(.A(G176gat), .B1(new_n933_), .B2(new_n633_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n881_), .A2(KEYINPUT124), .A3(new_n511_), .ZN(new_n935_));
  AOI21_X1  g734(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n511_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n925_), .A2(new_n212_), .A3(new_n632_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n934_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n927_), .A2(new_n280_), .A3(new_n674_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n925_), .A2(new_n674_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n935_), .B2(new_n936_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n942_), .B2(new_n204_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n927_), .B2(new_n742_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n753_), .A2(new_n203_), .A3(new_n209_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n927_), .B2(new_n945_), .ZN(G1351gat));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947_));
  NOR4_X1   g746(.A1(new_n537_), .A2(new_n461_), .A3(new_n511_), .A4(new_n350_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n881_), .A2(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n573_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n947_), .B1(new_n950_), .B2(G197gat), .ZN(new_n951_));
  OAI211_X1 g750(.A(KEYINPUT125), .B(new_n256_), .C1(new_n949_), .C2(new_n573_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(G197gat), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(G1352gat));
  NOR2_X1   g753(.A1(new_n949_), .A2(new_n632_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(new_n254_), .ZN(G1353gat));
  NOR2_X1   g755(.A1(new_n949_), .A2(new_n674_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(KEYINPUT126), .B1(new_n957_), .B2(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961_));
  OAI211_X1 g760(.A(new_n961_), .B(new_n958_), .C1(new_n949_), .C2(new_n674_), .ZN(new_n962_));
  XOR2_X1   g761(.A(KEYINPUT63), .B(G211gat), .Z(new_n963_));
  AOI22_X1  g762(.A1(new_n960_), .A2(new_n962_), .B1(new_n957_), .B2(new_n963_), .ZN(G1354gat));
  INV_X1    g763(.A(new_n949_), .ZN(new_n965_));
  AOI21_X1  g764(.A(G218gat), .B1(new_n965_), .B2(new_n753_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n704_), .A2(G218gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT127), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n965_), .B2(new_n968_), .ZN(G1355gat));
endmodule


