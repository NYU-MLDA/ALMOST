//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205_));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(G29gat), .B(G36gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G29gat), .B(G36gat), .Z(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n205_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(new_n211_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n212_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT15), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n225_), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(KEYINPUT64), .A3(new_n227_), .A4(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  AND3_X1   g029(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(KEYINPUT65), .A3(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT9), .ZN(new_n241_));
  AND2_X1   g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G85gat), .A2(G92gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n241_), .B1(new_n244_), .B2(KEYINPUT9), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n229_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n248_));
  INV_X1    g047(.A(G85gat), .ZN(new_n249_));
  INV_X1    g048(.A(G92gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(KEYINPUT67), .A3(new_n240_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT8), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT7), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT66), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n261_), .A3(new_n258_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n256_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n254_), .B1(new_n239_), .B2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n231_), .A2(new_n232_), .ZN(new_n265_));
  NOR4_X1   g064(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n261_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n265_), .B(new_n255_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n248_), .A2(new_n252_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n253_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n246_), .B1(new_n264_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n221_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n204_), .B1(new_n272_), .B2(KEYINPUT73), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n236_), .A2(new_n237_), .A3(new_n255_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n248_), .A2(new_n252_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT8), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n255_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n233_), .A2(new_n238_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n253_), .B(new_n269_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n213_), .A2(new_n214_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n246_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n272_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n274_), .A2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n272_), .A2(new_n284_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n273_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G134gat), .B(G162gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT36), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n290_), .A2(new_n297_), .A3(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT37), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n286_), .A2(new_n289_), .A3(KEYINPUT36), .A4(new_n296_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n301_), .A2(KEYINPUT76), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n297_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n298_), .B(new_n291_), .C1(new_n286_), .C2(new_n289_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n303_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n302_), .A2(KEYINPUT76), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(KEYINPUT76), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(G1gat), .ZN(new_n313_));
  INV_X1    g112(.A(G8gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT14), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G8gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G231gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G57gat), .B(G64gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT11), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT11), .ZN(new_n324_));
  INV_X1    g123(.A(G57gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(G64gat), .ZN(new_n326_));
  INV_X1    g125(.A(G64gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(G57gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n324_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(G71gat), .A2(G78gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G71gat), .A2(G78gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n323_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(G57gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(G64gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT11), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G71gat), .B(G78gat), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n336_), .A2(KEYINPUT68), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n322_), .B1(new_n333_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT68), .B1(new_n336_), .B2(new_n337_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n322_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n332_), .B(new_n323_), .C1(new_n321_), .C2(KEYINPUT11), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n320_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G183gat), .B(G211gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT17), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(KEYINPUT17), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n345_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n345_), .A2(new_n351_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n311_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G230gat), .ZN(new_n358_));
  INV_X1    g157(.A(G233gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n341_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n271_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n344_), .A2(new_n282_), .A3(new_n246_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n361_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT12), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT12), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n271_), .A2(new_n371_), .A3(new_n364_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n361_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G120gat), .B(G148gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G204gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT5), .B(G176gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT70), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n369_), .A2(new_n379_), .A3(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT13), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n357_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT78), .Z(new_n387_));
  INV_X1    g186(.A(KEYINPUT95), .ZN(new_n388_));
  XOR2_X1   g187(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  OR2_X1    g192(.A1(G197gat), .A2(G204gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT88), .B(G204gat), .Z(new_n395_));
  INV_X1    g194(.A(G197gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT89), .ZN(new_n398_));
  XOR2_X1   g197(.A(G211gat), .B(G218gat), .Z(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT21), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT21), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(new_n396_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(G197gat), .B2(G204gat), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n402_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT22), .B(G169gat), .ZN(new_n408_));
  INV_X1    g207(.A(G176gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G183gat), .ZN(new_n414_));
  INV_X1    g213(.A(G190gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT81), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT23), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G183gat), .A2(G190gat), .ZN(new_n418_));
  OAI22_X1  g217(.A1(new_n413_), .A2(KEYINPUT93), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n413_), .A2(KEYINPUT93), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT25), .B(G183gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(G190gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(G169gat), .A2(G176gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(KEYINPUT24), .A3(new_n411_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n423_), .B(new_n425_), .C1(KEYINPUT24), .C2(new_n424_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT23), .Z(new_n428_));
  OAI22_X1  g227(.A1(new_n419_), .A2(new_n420_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n407_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT22), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n409_), .B1(new_n431_), .B2(KEYINPUT82), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G169gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n432_), .A2(G169gat), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n433_), .B(new_n434_), .C1(new_n428_), .C2(new_n418_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n417_), .B2(new_n426_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n407_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT19), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n430_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n439_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n440_), .B1(new_n407_), .B2(new_n429_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n426_), .A2(new_n417_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n400_), .A2(new_n406_), .A3(new_n445_), .A4(new_n435_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n393_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n439_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n393_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n430_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n388_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n448_), .A2(new_n453_), .A3(new_n388_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT98), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT84), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464_));
  AND2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n464_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n459_), .B(new_n461_), .C1(new_n466_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n465_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n459_), .A2(KEYINPUT87), .ZN(new_n472_));
  AOI22_X1  g271(.A1(KEYINPUT3), .A2(new_n461_), .B1(new_n472_), .B2(KEYINPUT2), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(KEYINPUT2), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT86), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n463_), .B(new_n471_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n470_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G127gat), .B(G134gat), .Z(new_n480_));
  XOR2_X1   g279(.A(G113gat), .B(G120gat), .Z(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n470_), .A3(new_n478_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G225gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT96), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(KEYINPUT4), .A3(new_n485_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT4), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n479_), .A2(new_n491_), .A3(new_n482_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n488_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G29gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT0), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(new_n325_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G85gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT97), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(KEYINPUT33), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n495_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n499_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n457_), .A2(new_n458_), .A3(new_n503_), .A4(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n448_), .A2(new_n453_), .A3(new_n388_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n508_), .B(new_n503_), .C1(new_n510_), .C2(new_n454_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT98), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n495_), .A2(new_n499_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT100), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT100), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n500_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n449_), .A2(new_n439_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT99), .B(KEYINPUT20), .Z(new_n518_));
  NAND3_X1  g317(.A1(new_n430_), .A2(new_n437_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n439_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n450_), .A2(new_n452_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n451_), .A2(KEYINPUT32), .ZN(new_n522_));
  MUX2_X1   g321(.A(new_n520_), .B(new_n521_), .S(new_n522_), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n509_), .A2(new_n512_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n436_), .B(KEYINPUT30), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT83), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT31), .ZN(new_n528_));
  XOR2_X1   g327(.A(G71gat), .B(G99gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G43gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G227gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n484_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n527_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n479_), .A2(KEYINPUT29), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n407_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G228gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n359_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n407_), .B(new_n542_), .C1(new_n544_), .C2(new_n359_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G78gat), .B(G106gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n547_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n548_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n546_), .A2(KEYINPUT91), .A3(new_n547_), .A4(new_n549_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n479_), .A2(KEYINPUT29), .ZN(new_n556_));
  XOR2_X1   g355(.A(G22gat), .B(G50gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT28), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n556_), .B(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n554_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(new_n559_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n554_), .A2(new_n563_), .A3(new_n550_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n541_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n525_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n516_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT27), .B(new_n453_), .C1(new_n520_), .C2(new_n451_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT27), .ZN(new_n573_));
  INV_X1    g372(.A(new_n453_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n451_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n562_), .A2(new_n567_), .A3(new_n540_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n540_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n571_), .B(new_n577_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n570_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n318_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n215_), .B2(new_n220_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n283_), .A2(new_n582_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n318_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n318_), .B(KEYINPUT79), .C1(new_n213_), .C2(new_n214_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n585_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT80), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n594_), .B(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n387_), .A2(new_n581_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n313_), .A3(new_n516_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n307_), .B1(new_n570_), .B2(new_n580_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(new_n385_), .A3(new_n355_), .A4(new_n600_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n571_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n603_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT101), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT40), .ZN(new_n611_));
  OAI21_X1  g410(.A(G8gat), .B1(new_n606_), .B2(new_n577_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT102), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT102), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n612_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n577_), .A2(G8gat), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n601_), .A2(new_n617_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT103), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(KEYINPUT103), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n611_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT40), .A3(new_n620_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(G1325gat));
  OAI21_X1  g425(.A(G15gat), .B1(new_n606_), .B2(new_n541_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT41), .Z(new_n628_));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n601_), .A2(new_n629_), .A3(new_n540_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1326gat));
  NAND2_X1  g430(.A1(new_n562_), .A2(new_n567_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n606_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n601_), .A2(new_n636_), .A3(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1327gat));
  NAND2_X1  g437(.A1(new_n385_), .A2(new_n600_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n355_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n581_), .A2(new_n307_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT107), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT107), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n581_), .A2(new_n640_), .A3(new_n643_), .A4(new_n307_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n516_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  INV_X1    g446(.A(new_n311_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n648_), .B1(new_n570_), .B2(new_n580_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n571_), .A2(new_n577_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n579_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n562_), .A2(new_n567_), .A3(new_n540_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n511_), .A2(KEYINPUT98), .B1(new_n516_), .B2(new_n523_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n568_), .B1(new_n656_), .B2(new_n509_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n311_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n650_), .B(new_n311_), .C1(new_n655_), .C2(new_n657_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n651_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n640_), .B(KEYINPUT104), .Z(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT106), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n666_), .B(KEYINPUT44), .C1(new_n661_), .C2(new_n662_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n662_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n670_), .A2(G29gat), .A3(new_n516_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n646_), .B1(new_n669_), .B2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(KEYINPUT108), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n577_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n670_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n577_), .A2(G36gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n642_), .A2(new_n644_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT45), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n642_), .A2(new_n644_), .A3(new_n682_), .A4(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n673_), .A2(KEYINPUT108), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n675_), .B1(new_n678_), .B2(new_n687_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n674_), .B(new_n686_), .C1(new_n677_), .C2(G36gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  AOI21_X1  g489(.A(G43gat), .B1(new_n645_), .B2(new_n540_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n670_), .A2(G43gat), .A3(new_n540_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n668_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g494(.A(G50gat), .B1(new_n645_), .B2(new_n632_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n670_), .A2(G50gat), .A3(new_n632_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n669_), .B2(new_n697_), .ZN(G1331gat));
  INV_X1    g497(.A(new_n600_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n384_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n581_), .A2(new_n357_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n325_), .A3(new_n516_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n605_), .A2(new_n355_), .A3(new_n701_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G57gat), .B1(new_n705_), .B2(new_n571_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1332gat));
  OAI21_X1  g506(.A(G64gat), .B1(new_n705_), .B2(new_n577_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT109), .Z(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n703_), .A2(new_n327_), .A3(new_n676_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1333gat));
  OAI21_X1  g511(.A(G71gat), .B1(new_n705_), .B2(new_n541_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n541_), .A2(G71gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n702_), .B2(new_n716_), .ZN(G1334gat));
  OAI21_X1  g516(.A(G78gat), .B1(new_n705_), .B2(new_n633_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT111), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n702_), .A2(G78gat), .A3(new_n633_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1335gat));
  NOR2_X1   g521(.A1(new_n700_), .A2(new_n355_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n581_), .A2(new_n307_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n249_), .A3(new_n516_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n723_), .B(KEYINPUT112), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT105), .B1(new_n658_), .B2(KEYINPUT43), .ZN(new_n728_));
  INV_X1    g527(.A(new_n660_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n730_), .B2(new_n659_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n516_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n726_), .B1(new_n732_), .B2(new_n249_), .ZN(G1336gat));
  NAND3_X1  g532(.A1(new_n725_), .A2(new_n250_), .A3(new_n676_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n731_), .A2(new_n676_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n250_), .ZN(G1337gat));
  NOR3_X1   g535(.A1(new_n724_), .A2(new_n225_), .A3(new_n541_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n731_), .A2(new_n540_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G99gat), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT51), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n739_), .B(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n227_), .A3(new_n632_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n731_), .A2(new_n632_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(G106gat), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT52), .B(new_n227_), .C1(new_n731_), .C2(new_n632_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g548(.A1(new_n676_), .A2(new_n571_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n578_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(KEYINPUT59), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT54), .B1(new_n386_), .B2(new_n600_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n357_), .A2(new_n755_), .A3(new_n385_), .A4(new_n699_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n307_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n600_), .A2(new_n382_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n360_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n361_), .A2(KEYINPUT114), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(KEYINPUT55), .A2(new_n761_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n763_), .A2(new_n765_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n380_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  OAI211_X1 g569(.A(KEYINPUT56), .B(new_n380_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n760_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n584_), .A2(KEYINPUT115), .A3(new_n586_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT115), .ZN(new_n774_));
  INV_X1    g573(.A(new_n586_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n583_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n592_), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n590_), .A2(new_n591_), .A3(new_n585_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n598_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n594_), .A2(new_n599_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n383_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n759_), .B1(new_n772_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT57), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n382_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n771_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n374_), .A2(new_n762_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n373_), .A2(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n764_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n763_), .A2(new_n765_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n380_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT58), .B(new_n785_), .C1(new_n786_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n784_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT58), .B1(new_n796_), .B2(KEYINPUT116), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n785_), .B1(new_n786_), .B2(new_n792_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n797_), .A2(new_n800_), .B1(new_n310_), .B2(new_n304_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n795_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n796_), .A2(KEYINPUT116), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n311_), .B(new_n802_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n783_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n356_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n758_), .B1(new_n810_), .B2(KEYINPUT121), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n810_), .A2(KEYINPUT121), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n753_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(G113gat), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(G113gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n600_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n783_), .B(KEYINPUT119), .C1(new_n803_), .C2(new_n808_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n356_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n751_), .B1(new_n821_), .B2(new_n757_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT120), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n355_), .B1(new_n809_), .B2(new_n818_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n758_), .B1(new_n826_), .B2(new_n820_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(KEYINPUT59), .C1(new_n827_), .C2(new_n751_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n813_), .B(new_n817_), .C1(new_n824_), .C2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G113gat), .B1(new_n822_), .B2(new_n600_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT123), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n824_), .A2(new_n828_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n813_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n817_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  INV_X1    g635(.A(new_n830_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(G1340gat));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  AOI21_X1  g639(.A(G120gat), .B1(new_n384_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(G120gat), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n841_), .A2(new_n842_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n822_), .A2(new_n843_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n813_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n847_), .A2(new_n384_), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n846_), .B1(new_n848_), .B2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n822_), .B2(new_n355_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT125), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n355_), .A2(G127gat), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(KEYINPUT126), .Z(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n847_), .B2(new_n854_), .ZN(G1342gat));
  INV_X1    g654(.A(G134gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n822_), .A2(new_n856_), .A3(new_n307_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n847_), .A2(new_n311_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n827_), .A2(new_n653_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n750_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n699_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n385_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT127), .B(G148gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NOR2_X1   g665(.A1(new_n861_), .A2(new_n356_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT61), .B(G155gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n861_), .B2(new_n648_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n759_), .A2(G162gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n861_), .B2(new_n871_), .ZN(G1347gat));
  NAND2_X1  g671(.A1(new_n811_), .A2(new_n812_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n577_), .A2(new_n516_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n540_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n632_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877_), .B2(new_n699_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n877_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n408_), .A3(new_n600_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n879_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n882_), .A3(new_n883_), .ZN(G1348gat));
  AOI21_X1  g683(.A(G176gat), .B1(new_n881_), .B2(new_n384_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n827_), .A2(new_n632_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n875_), .A2(new_n385_), .A3(new_n409_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  NOR3_X1   g687(.A1(new_n877_), .A2(new_n356_), .A3(new_n421_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n886_), .A2(new_n355_), .A3(new_n540_), .A4(new_n874_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n414_), .B2(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n877_), .B2(new_n648_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n307_), .A2(new_n422_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n877_), .B2(new_n893_), .ZN(G1351gat));
  NAND2_X1  g693(.A1(new_n860_), .A2(new_n874_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n699_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n396_), .ZN(G1352gat));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n385_), .ZN(new_n898_));
  MUX2_X1   g697(.A(G204gat), .B(new_n395_), .S(new_n898_), .Z(G1353gat));
  NAND3_X1  g698(.A1(new_n860_), .A2(new_n355_), .A3(new_n874_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  OAI21_X1  g703(.A(G218gat), .B1(new_n895_), .B2(new_n648_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n759_), .A2(G218gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n895_), .B2(new_n906_), .ZN(G1355gat));
endmodule


