//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n206_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n206_), .C1(new_n211_), .C2(new_n217_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n223_), .B1(new_n226_), .B2(new_n214_), .ZN(new_n227_));
  NOR4_X1   g026(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT64), .A4(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n208_), .A2(new_n210_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT9), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n205_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n204_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n231_), .B1(new_n205_), .B2(new_n232_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n230_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n229_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT10), .B(G99gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT64), .B1(new_n239_), .B2(G106gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n226_), .A2(new_n223_), .A3(new_n214_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n205_), .A2(new_n232_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT65), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n245_), .A2(new_n233_), .A3(new_n204_), .A4(new_n234_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n242_), .A2(new_n243_), .A3(new_n246_), .A4(new_n230_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n222_), .A2(new_n238_), .A3(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n248_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT73), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n246_), .B(new_n230_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(KEYINPUT66), .A2(new_n258_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(new_n253_), .A3(new_n247_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT35), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n257_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n263_), .A2(new_n264_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n256_), .A2(KEYINPUT73), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT74), .ZN(new_n272_));
  XOR2_X1   g071(.A(G134gat), .B(G162gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT36), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n267_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n270_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n274_), .B(KEYINPUT36), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(KEYINPUT11), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n286_));
  XOR2_X1   g085(.A(G71gat), .B(G78gat), .Z(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n282_), .A3(KEYINPUT11), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(KEYINPUT11), .B2(new_n283_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(new_n284_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n293_), .B1(new_n259_), .B2(new_n247_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n293_), .A2(new_n222_), .A3(new_n238_), .A4(new_n247_), .ZN(new_n300_));
  INV_X1    g099(.A(G230gat), .ZN(new_n301_));
  INV_X1    g100(.A(G233gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT69), .B1(new_n299_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n248_), .A2(new_n294_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n297_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .A4(new_n295_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n300_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n303_), .B1(new_n313_), .B2(new_n296_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT5), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G176gat), .B(G204gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n314_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(KEYINPUT70), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n315_), .A2(new_n324_), .A3(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT13), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(KEYINPUT13), .A3(new_n325_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(KEYINPUT71), .A3(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G15gat), .B(G22gat), .ZN(new_n336_));
  INV_X1    g135(.A(G1gat), .ZN(new_n337_));
  INV_X1    g136(.A(G8gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT14), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G8gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n255_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n253_), .A3(new_n343_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G229gat), .A2(G233gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n344_), .B(new_n253_), .Z(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G229gat), .A3(G233gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G113gat), .B(G141gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT78), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G169gat), .B(G197gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n349_), .A2(new_n351_), .A3(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n335_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G231gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n344_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(new_n293_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT17), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G127gat), .B(G155gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT16), .ZN(new_n367_));
  XOR2_X1   g166(.A(G183gat), .B(G211gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n364_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(KEYINPUT17), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n364_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G15gat), .B(G43gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT80), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT30), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT23), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(G183gat), .B2(G190gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G169gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(KEYINPUT24), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT79), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT25), .B(G183gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n384_), .A2(KEYINPUT24), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n377_), .A3(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n381_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n375_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(G71gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n394_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G127gat), .B(G134gat), .Z(new_n400_));
  XOR2_X1   g199(.A(G113gat), .B(G120gat), .Z(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n400_), .A2(new_n401_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n404_), .B2(new_n403_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT31), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(new_n213_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n399_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n399_), .A2(new_n408_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G22gat), .B(G50gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G141gat), .A2(G148gat), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n414_), .A2(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n415_), .B2(new_n414_), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n417_), .B(KEYINPUT82), .Z(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G155gat), .A2(G162gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT83), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G155gat), .A3(G162gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G155gat), .ZN(new_n428_));
  INV_X1    g227(.A(G162gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n422_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n430_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n434_));
  OAI221_X1 g233(.A(new_n420_), .B1(G141gat), .B2(G148gat), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT85), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n431_), .A2(new_n438_), .A3(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT29), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n413_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n413_), .A3(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n437_), .A2(KEYINPUT29), .A3(new_n439_), .ZN(new_n451_));
  AND2_X1   g250(.A1(G228gat), .A2(G233gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G211gat), .B(G218gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(G197gat), .B(G204gat), .Z(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(KEYINPUT87), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(KEYINPUT21), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n455_), .B(KEYINPUT21), .C1(new_n454_), .C2(new_n453_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n452_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n436_), .A2(KEYINPUT29), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n457_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n451_), .A2(new_n458_), .B1(new_n461_), .B2(new_n452_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n464_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n450_), .A2(KEYINPUT88), .A3(new_n465_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n449_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n462_), .A2(new_n464_), .ZN(new_n469_));
  OAI22_X1  g268(.A1(new_n468_), .A2(new_n447_), .B1(KEYINPUT88), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n467_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n437_), .A2(new_n406_), .A3(new_n439_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n403_), .A2(new_n402_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n431_), .A2(new_n435_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT94), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n431_), .A2(new_n435_), .A3(new_n478_), .A4(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G85gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT0), .B(G57gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  AND3_X1   g285(.A1(new_n474_), .A2(new_n480_), .A3(KEYINPUT4), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n481_), .B(KEYINPUT95), .Z(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n474_), .B2(KEYINPUT4), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n482_), .B(new_n486_), .C1(new_n487_), .C2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT96), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n474_), .A2(new_n480_), .A3(KEYINPUT4), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n488_), .C1(KEYINPUT4), .C2(new_n474_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n494_), .A2(KEYINPUT96), .A3(new_n482_), .A4(new_n486_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT33), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT97), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n385_), .A2(KEYINPUT24), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n499_), .A2(new_n500_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n385_), .A2(KEYINPUT89), .A3(KEYINPUT24), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n381_), .B1(new_n503_), .B2(new_n392_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n460_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G226gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT19), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT90), .B1(new_n460_), .B2(new_n393_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n460_), .A2(KEYINPUT90), .A3(new_n393_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n507_), .B(new_n510_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n460_), .A2(new_n504_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(KEYINPUT20), .C1(new_n393_), .C2(new_n460_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n509_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G8gat), .B(G36gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(G64gat), .B(G92gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT92), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT93), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n513_), .A2(new_n516_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n521_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI211_X1 g328(.A(KEYINPUT93), .B(new_n521_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n524_), .B(new_n525_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n486_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n474_), .A2(new_n480_), .A3(new_n488_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n481_), .B1(new_n474_), .B2(KEYINPUT4), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n533_), .C1(new_n487_), .C2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n490_), .B2(new_n496_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n492_), .A2(new_n495_), .A3(new_n538_), .A4(new_n496_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n498_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n494_), .A2(new_n482_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n532_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n490_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n507_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n509_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n521_), .A2(KEYINPUT32), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT98), .B1(new_n527_), .B2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT98), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n543_), .B(new_n550_), .C1(new_n551_), .C2(new_n548_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n473_), .B1(new_n540_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n543_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n472_), .A3(new_n467_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT27), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n531_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n546_), .A2(new_n528_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT27), .A3(new_n522_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n411_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n473_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n560_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n411_), .A2(new_n543_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  AND4_X1   g366(.A1(new_n281_), .A2(new_n361_), .A3(new_n372_), .A4(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n543_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G1gat), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT38), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n562_), .A2(new_n566_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n360_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  OAI211_X1 g374(.A(KEYINPUT75), .B(new_n575_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n278_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n276_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n578_), .B2(new_n269_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n270_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n575_), .A2(KEYINPUT75), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n575_), .A2(KEYINPUT75), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n576_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n372_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n574_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n576_), .A2(KEYINPUT76), .A3(new_n583_), .A4(new_n372_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n334_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n573_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n572_), .B(new_n591_), .C1(new_n590_), .C2(new_n589_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n337_), .A3(new_n543_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n593_), .A2(KEYINPUT99), .A3(new_n571_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT99), .B1(new_n593_), .B2(new_n571_), .ZN(new_n595_));
  OAI221_X1 g394(.A(new_n570_), .B1(new_n571_), .B2(new_n593_), .C1(new_n594_), .C2(new_n595_), .ZN(G1324gat));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n338_), .A3(new_n560_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n568_), .A2(new_n560_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(G8gat), .ZN(new_n600_));
  AOI211_X1 g399(.A(KEYINPUT39), .B(new_n338_), .C1(new_n568_), .C2(new_n560_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g402(.A(G15gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n411_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n592_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n568_), .A2(new_n605_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n608_));
  AND3_X1   g407(.A1(new_n607_), .A2(G15gat), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n607_), .B2(G15gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n606_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(G1326gat));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n592_), .A2(new_n614_), .A3(new_n473_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n568_), .A2(new_n473_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(G22gat), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(KEYINPUT42), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(KEYINPUT42), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(G1327gat));
  NOR2_X1   g419(.A1(new_n281_), .A2(new_n372_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n361_), .A2(new_n567_), .A3(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n554_), .A2(G29gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT104), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n335_), .A2(new_n360_), .A3(new_n372_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n567_), .B2(new_n584_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n584_), .ZN(new_n629_));
  AOI211_X1 g428(.A(KEYINPUT43), .B(new_n629_), .C1(new_n562_), .C2(new_n566_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT44), .B(new_n626_), .C1(new_n628_), .C2(new_n630_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n543_), .A4(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n543_), .A3(new_n635_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT102), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n637_), .A2(KEYINPUT103), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT103), .B1(new_n637_), .B2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n625_), .B1(new_n640_), .B2(new_n641_), .ZN(G1328gat));
  NOR2_X1   g441(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT46), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n647_), .A3(new_n560_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n633_), .A2(new_n560_), .A3(new_n635_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G36gat), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n643_), .B(new_n646_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n652_));
  AND4_X1   g451(.A1(new_n644_), .A2(new_n649_), .A3(new_n645_), .A4(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND3_X1  g453(.A1(new_n633_), .A2(new_n605_), .A3(new_n635_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G43gat), .ZN(new_n656_));
  INV_X1    g455(.A(G43gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n622_), .A2(new_n657_), .A3(new_n605_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1330gat));
  AOI21_X1  g460(.A(G50gat), .B1(new_n622_), .B2(new_n473_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n633_), .A2(new_n635_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n473_), .A2(G50gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(G1331gat));
  NAND3_X1  g464(.A1(new_n335_), .A2(new_n360_), .A3(new_n372_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n666_), .A2(new_n572_), .A3(new_n280_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(G57gat), .A3(new_n543_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT111), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n588_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT107), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n588_), .A2(new_n332_), .A3(new_n672_), .A4(new_n333_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n567_), .B2(new_n360_), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT108), .B(new_n573_), .C1(new_n562_), .C2(new_n566_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT109), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n674_), .B(new_n680_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n679_), .A2(KEYINPUT110), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT110), .B1(new_n679_), .B2(new_n681_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n554_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n669_), .B1(new_n684_), .B2(G57gat), .ZN(new_n685_));
  INV_X1    g484(.A(G57gat), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n678_), .A2(KEYINPUT109), .ZN(new_n688_));
  INV_X1    g487(.A(new_n681_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n543_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT111), .B(new_n686_), .C1(new_n691_), .C2(new_n682_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n668_), .B1(new_n685_), .B2(new_n692_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n667_), .B2(new_n560_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT48), .Z(new_n696_));
  NOR2_X1   g495(.A1(new_n688_), .A2(new_n689_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(new_n694_), .A3(new_n560_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1333gat));
  AOI21_X1  g498(.A(new_n396_), .B1(new_n667_), .B2(new_n605_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT49), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n396_), .A3(new_n605_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1334gat));
  INV_X1    g502(.A(G78gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n667_), .B2(new_n473_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT50), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n704_), .A3(new_n473_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1335gat));
  NOR2_X1   g507(.A1(new_n676_), .A2(new_n677_), .ZN(new_n709_));
  NOR4_X1   g508(.A1(new_n709_), .A2(new_n281_), .A3(new_n372_), .A4(new_n334_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n202_), .A3(new_n543_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n335_), .A2(new_n360_), .A3(new_n585_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT112), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n628_), .A2(new_n630_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n543_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n716_), .B2(new_n202_), .ZN(G1336gat));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n560_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n564_), .A2(G92gat), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n718_), .A2(G92gat), .B1(new_n710_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1337gat));
  NAND2_X1  g521(.A1(new_n715_), .A2(new_n605_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n411_), .A2(new_n239_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n723_), .A2(G99gat), .B1(new_n710_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1338gat));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n214_), .A3(new_n473_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n473_), .A3(new_n714_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(new_n728_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  NAND4_X1  g536(.A1(new_n330_), .A2(new_n360_), .A3(new_n629_), .A4(new_n372_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT54), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n573_), .A2(new_n322_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n306_), .A2(new_n741_), .A3(new_n311_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT114), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n306_), .A2(new_n744_), .A3(new_n741_), .A4(new_n311_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n303_), .B1(new_n299_), .B2(new_n313_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT55), .A4(new_n295_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AND4_X1   g548(.A1(KEYINPUT115), .A2(new_n743_), .A3(new_n745_), .A4(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n742_), .B2(KEYINPUT114), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT115), .B1(new_n751_), .B2(new_n745_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n319_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n743_), .A2(new_n745_), .A3(new_n749_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n751_), .A2(KEYINPUT115), .A3(new_n745_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n319_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n740_), .B1(new_n755_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n358_), .B1(new_n350_), .B2(new_n348_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n347_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n348_), .ZN(new_n765_));
  AND4_X1   g564(.A1(new_n359_), .A2(new_n323_), .A3(new_n325_), .A4(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n281_), .B1(new_n762_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT57), .B(new_n281_), .C1(new_n762_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n755_), .A2(new_n761_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n322_), .A2(new_n359_), .A3(new_n765_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT58), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n319_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n754_), .B(new_n321_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT58), .B(new_n772_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n584_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n769_), .B(new_n770_), .C1(new_n773_), .C2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n739_), .B1(new_n778_), .B2(new_n585_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n473_), .A2(new_n560_), .A3(new_n411_), .A4(new_n554_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OR3_X1    g581(.A1(new_n779_), .A2(KEYINPUT118), .A3(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT118), .B1(new_n779_), .B2(new_n782_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n777_), .B2(new_n773_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n772_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n789_), .A2(KEYINPUT117), .A3(new_n584_), .A4(new_n776_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n770_), .A4(new_n769_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n585_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n739_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n780_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n783_), .B(new_n784_), .C1(new_n781_), .C2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G113gat), .B1(new_n797_), .B2(new_n360_), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n795_), .A2(G113gat), .A3(new_n360_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1340gat));
  OAI21_X1  g599(.A(G120gat), .B1(new_n797_), .B2(new_n334_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT60), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT119), .B1(new_n802_), .B2(G120gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(G120gat), .B1(new_n335_), .B2(new_n802_), .ZN(new_n804_));
  MUX2_X1   g603(.A(new_n803_), .B(KEYINPUT119), .S(new_n804_), .Z(new_n805_));
  NAND2_X1  g604(.A1(new_n796_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n801_), .A2(new_n806_), .ZN(G1341gat));
  OAI21_X1  g606(.A(G127gat), .B1(new_n797_), .B2(new_n585_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n795_), .A2(G127gat), .A3(new_n585_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1342gat));
  OAI21_X1  g609(.A(G134gat), .B1(new_n797_), .B2(new_n629_), .ZN(new_n811_));
  OR3_X1    g610(.A1(new_n795_), .A2(G134gat), .A3(new_n281_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(G1343gat));
  NOR4_X1   g612(.A1(new_n563_), .A2(new_n605_), .A3(new_n554_), .A4(new_n560_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n573_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n335_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n372_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT61), .B(G155gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1346gat));
  NAND3_X1  g622(.A1(new_n816_), .A2(G162gat), .A3(new_n584_), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT120), .B(G162gat), .C1(new_n816_), .C2(new_n280_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n794_), .A2(new_n280_), .A3(new_n814_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n429_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT121), .B(new_n824_), .C1(new_n825_), .C2(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1347gat));
  NAND2_X1  g632(.A1(new_n565_), .A2(new_n560_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n779_), .A2(new_n473_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT22), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n573_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G169gat), .ZN(new_n841_));
  INV_X1    g640(.A(new_n835_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n360_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n382_), .B1(new_n843_), .B2(new_n838_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n844_), .B2(new_n840_), .ZN(G1348gat));
  OAI21_X1  g644(.A(new_n383_), .B1(new_n842_), .B2(new_n334_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n794_), .A2(KEYINPUT123), .A3(new_n563_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n739_), .B1(new_n791_), .B2(new_n585_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n473_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n834_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n334_), .A2(new_n383_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n847_), .A2(new_n850_), .A3(new_n851_), .A4(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n846_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n846_), .A2(KEYINPUT124), .A3(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1349gat));
  NOR3_X1   g657(.A1(new_n842_), .A2(new_n585_), .A3(new_n388_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n847_), .A2(new_n850_), .A3(new_n372_), .A4(new_n851_), .ZN(new_n860_));
  INV_X1    g659(.A(G183gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n842_), .B2(new_n629_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n835_), .A2(new_n280_), .A3(new_n389_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1351gat));
  NOR3_X1   g664(.A1(new_n555_), .A2(new_n564_), .A3(new_n605_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n794_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n573_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n794_), .A2(new_n866_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n334_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT125), .B(G204gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1353gat));
  NAND2_X1  g672(.A1(new_n867_), .A2(new_n372_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT63), .B(G211gat), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n877_));
  INV_X1    g676(.A(G211gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n874_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n874_), .A2(KEYINPUT126), .A3(new_n877_), .A4(new_n878_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n876_), .B1(new_n881_), .B2(new_n882_), .ZN(G1354gat));
  AND3_X1   g682(.A1(new_n867_), .A2(G218gat), .A3(new_n584_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n870_), .A2(KEYINPUT127), .A3(new_n281_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(G218gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT127), .B1(new_n870_), .B2(new_n281_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(G1355gat));
endmodule


