//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT82), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT23), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G190gat), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n211_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT26), .B1(new_n211_), .B2(KEYINPUT81), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n208_), .B(new_n210_), .C1(new_n212_), .C2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT30), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G71gat), .B(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n221_), .B(KEYINPUT30), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n224_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT83), .B(G43gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT84), .B(G15gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT86), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n226_), .A2(new_n228_), .A3(new_n234_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G113gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G120gat), .ZN(new_n246_));
  INV_X1    g045(.A(G113gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n244_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G120gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT31), .Z(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n236_), .A2(KEYINPUT87), .A3(new_n238_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n241_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n239_), .A2(new_n240_), .A3(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259_));
  INV_X1    g058(.A(G141gat), .ZN(new_n260_));
  INV_X1    g059(.A(G148gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n262_), .A2(new_n265_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G155gat), .B(G162gat), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT88), .ZN(new_n271_));
  INV_X1    g070(.A(G155gat), .ZN(new_n272_));
  INV_X1    g071(.A(G162gat), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n272_), .A2(new_n273_), .A3(KEYINPUT1), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT1), .B1(new_n272_), .B2(new_n273_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n274_), .B(new_n275_), .C1(G155gat), .C2(G162gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n260_), .A2(new_n261_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n263_), .A3(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT92), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n251_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n251_), .A2(new_n280_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT4), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G225gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n279_), .A2(KEYINPUT4), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n251_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT93), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G1gat), .B(G29gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G85gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT0), .ZN(new_n292_));
  INV_X1    g091(.A(G57gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n283_), .A2(new_n296_), .A3(new_n285_), .A4(new_n287_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n289_), .A2(new_n294_), .A3(new_n295_), .A4(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT20), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT26), .B(G190gat), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n213_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n208_), .A2(new_n210_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT22), .B(G169gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT91), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n217_), .B(new_n209_), .C1(new_n307_), .C2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(G197gat), .B(G204gat), .Z(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(KEYINPUT21), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(KEYINPUT21), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  AOI21_X1  g113(.A(new_n301_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n221_), .B2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT19), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n309_), .A2(new_n314_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n221_), .A2(new_n314_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n318_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n320_), .A2(KEYINPUT20), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT18), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G64gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(G92gat), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n319_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n300_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n283_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n294_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n281_), .A2(new_n282_), .A3(new_n285_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n298_), .A2(KEYINPUT94), .A3(new_n299_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n298_), .A2(new_n299_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT94), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .A4(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n289_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n335_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n298_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n301_), .A2(KEYINPUT95), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n301_), .A2(KEYINPUT95), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n320_), .A2(new_n321_), .A3(new_n346_), .A4(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n318_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n318_), .B2(new_n316_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n328_), .A2(KEYINPUT32), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n345_), .B(new_n352_), .C1(new_n324_), .C2(new_n351_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n258_), .B1(new_n342_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G50gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n279_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT28), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(G22gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n358_), .A2(G22gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n355_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G50gat), .A3(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n314_), .B1(new_n279_), .B2(new_n356_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G78gat), .B(G106gat), .Z(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n369_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n373_), .A3(new_n371_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n365_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n370_), .A2(KEYINPUT90), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n370_), .A2(KEYINPUT90), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n375_), .B1(new_n378_), .B2(new_n365_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n354_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n350_), .A2(new_n329_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n331_), .A3(KEYINPUT27), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n332_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n257_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n362_), .A2(new_n364_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n388_), .A2(new_n373_), .A3(new_n377_), .A4(new_n376_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(new_n256_), .A3(new_n255_), .A4(new_n375_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n345_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n381_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G120gat), .B(G148gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT5), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G204gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(G85gat), .B(G92gat), .Z(new_n400_));
  NAND2_X1  g199(.A1(G99gat), .A2(G106gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G99gat), .A3(G106gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT7), .ZN(new_n406_));
  INV_X1    g205(.A(G99gat), .ZN(new_n407_));
  INV_X1    g206(.A(G106gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n400_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n403_), .B1(G99gat), .B2(G106gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n410_), .B(new_n409_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(KEYINPUT66), .A3(new_n400_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(KEYINPUT8), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT67), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G85gat), .B(G92gat), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n409_), .A2(new_n410_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n402_), .A2(new_n404_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT8), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n414_), .A2(new_n420_), .A3(KEYINPUT8), .A4(new_n418_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n400_), .A2(KEYINPUT9), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT64), .B(G92gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT9), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(G85gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n407_), .A2(KEYINPUT10), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n407_), .A2(KEYINPUT10), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n408_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n429_), .A2(new_n432_), .A3(new_n423_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT10), .B(G99gat), .Z(new_n439_));
  AOI22_X1  g238(.A1(new_n439_), .A2(new_n408_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n440_), .A2(KEYINPUT65), .A3(new_n429_), .A4(new_n432_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G78gat), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n445_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n427_), .A2(new_n428_), .A3(new_n442_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G230gat), .A2(G233gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT69), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n413_), .B(new_n421_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT66), .B1(new_n417_), .B2(new_n400_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n425_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n426_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n428_), .B(new_n442_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n449_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(KEYINPUT12), .A3(new_n449_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT69), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n451_), .A2(new_n464_), .A3(new_n452_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n454_), .A2(new_n462_), .A3(new_n463_), .A4(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT68), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n460_), .A2(new_n468_), .A3(new_n451_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n452_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n459_), .A2(KEYINPUT68), .A3(new_n449_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n467_), .B1(new_n466_), .B2(new_n472_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n399_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT13), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n466_), .A2(new_n472_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n480_), .A2(new_n399_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n478_), .B(new_n479_), .C1(new_n482_), .C2(new_n477_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n478_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n477_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT13), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT78), .B(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT14), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT79), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(G1gat), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT79), .ZN(new_n500_));
  INV_X1    g299(.A(G1gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(G8gat), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(G8gat), .B1(new_n498_), .B2(new_n502_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n504_), .A2(new_n505_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n498_), .A2(new_n502_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n491_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n514_), .B2(new_n503_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n489_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n489_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n510_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G113gat), .B(G141gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G169gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n522_), .B(G197gat), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n511_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n514_), .A2(new_n510_), .A3(new_n503_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n520_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n524_), .B1(new_n520_), .B2(new_n528_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n488_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n394_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n459_), .A2(new_n489_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n510_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT34), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT35), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n459_), .A2(new_n511_), .A3(new_n489_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(KEYINPUT35), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT72), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n535_), .A2(new_n538_), .A3(new_n539_), .A4(new_n542_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G134gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(new_n273_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n548_), .B(new_n552_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n547_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(KEYINPUT37), .B(new_n547_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n449_), .B(KEYINPUT80), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n514_), .A2(new_n503_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT16), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(G183gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(G211gat), .Z(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n566_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n561_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n533_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n345_), .A3(new_n490_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT38), .ZN(new_n581_));
  INV_X1    g380(.A(new_n556_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n533_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G1gat), .B1(new_n586_), .B2(new_n392_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n587_), .ZN(G1324gat));
  INV_X1    g387(.A(new_n386_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G8gat), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT97), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT97), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(KEYINPUT39), .A3(new_n592_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n579_), .A2(new_n491_), .A3(new_n386_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT96), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT40), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1325gat));
  INV_X1    g402(.A(G15gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n585_), .B2(new_n258_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT41), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n579_), .A2(new_n604_), .A3(new_n258_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  INV_X1    g407(.A(G22gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n585_), .B2(new_n379_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT42), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n579_), .A2(new_n609_), .A3(new_n379_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1327gat));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n394_), .B2(new_n561_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n354_), .A2(new_n380_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(KEYINPUT43), .A3(new_n560_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n532_), .B(new_n576_), .C1(new_n615_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT43), .B1(new_n616_), .B2(new_n560_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n394_), .A2(new_n614_), .A3(new_n561_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n623_), .A2(KEYINPUT44), .A3(new_n532_), .A4(new_n576_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(new_n345_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G29gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n532_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n616_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n582_), .A2(new_n583_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n392_), .A2(G29gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT98), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n626_), .B1(new_n630_), .B2(new_n632_), .ZN(G1328gat));
  INV_X1    g432(.A(KEYINPUT45), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n630_), .A2(G36gat), .A3(new_n589_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n635_), .A2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n636_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT45), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n642_), .A3(KEYINPUT101), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n620_), .A2(new_n386_), .A3(new_n624_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n620_), .A2(KEYINPUT99), .A3(new_n386_), .A4(new_n624_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(KEYINPUT101), .A3(G36gat), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n643_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1329gat));
  INV_X1    g451(.A(new_n630_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G43gat), .B1(new_n653_), .B2(new_n258_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT103), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n620_), .A2(G43gat), .A3(new_n258_), .A4(new_n624_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT47), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n655_), .B(new_n662_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1330gat));
  NAND3_X1  g463(.A1(new_n653_), .A2(new_n355_), .A3(new_n379_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n620_), .A2(new_n379_), .A3(new_n624_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G50gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G50gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1331gat));
  INV_X1    g469(.A(new_n531_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n487_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n394_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n584_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT105), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT106), .B1(new_n392_), .B2(new_n293_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n673_), .A2(new_n578_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n345_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n677_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n679_), .A2(new_n293_), .B1(new_n680_), .B2(KEYINPUT106), .ZN(G1332gat));
  INV_X1    g480(.A(G64gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n682_), .A3(new_n386_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n675_), .A2(new_n386_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G64gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT107), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(G64gat), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n686_), .A2(KEYINPUT48), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT48), .B1(new_n686_), .B2(new_n688_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n683_), .B1(new_n689_), .B2(new_n690_), .ZN(G1333gat));
  INV_X1    g490(.A(G71gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n678_), .A2(new_n692_), .A3(new_n258_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n675_), .B2(new_n258_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(new_n695_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT108), .B(new_n693_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1334gat));
  INV_X1    g501(.A(G78gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n675_), .B2(new_n379_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT50), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n678_), .A2(new_n703_), .A3(new_n379_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1335gat));
  NOR3_X1   g506(.A1(new_n673_), .A2(new_n583_), .A3(new_n582_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G85gat), .B1(new_n708_), .B2(new_n345_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n623_), .A2(new_n576_), .A3(new_n672_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n345_), .A2(G85gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(G1336gat));
  AOI21_X1  g511(.A(G92gat), .B1(new_n708_), .B2(new_n386_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n386_), .A2(new_n430_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n710_), .B2(new_n714_), .ZN(G1337gat));
  AOI21_X1  g514(.A(new_n407_), .B1(new_n710_), .B2(new_n258_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n258_), .A2(new_n439_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n708_), .B2(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g518(.A1(new_n708_), .A2(new_n408_), .A3(new_n379_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n710_), .A2(new_n379_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G106gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT52), .B(new_n408_), .C1(new_n710_), .C2(new_n379_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n459_), .A2(KEYINPUT12), .A3(new_n449_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT12), .B1(new_n459_), .B2(new_n449_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n451_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n731_), .B2(new_n452_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n466_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n462_), .A2(new_n463_), .A3(new_n451_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(KEYINPUT109), .A3(new_n470_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n728_), .A2(new_n729_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT55), .A3(new_n454_), .A4(new_n465_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n732_), .A2(new_n734_), .A3(new_n736_), .A4(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n399_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT56), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n399_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT56), .B1(new_n739_), .B2(new_n399_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n531_), .B1(new_n746_), .B2(KEYINPUT110), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n481_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n517_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n523_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT111), .B1(new_n750_), .B2(new_n524_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n518_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n519_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT112), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n516_), .A2(new_n759_), .A3(new_n519_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n760_), .A3(new_n749_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n529_), .B1(new_n755_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n748_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n582_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT58), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(KEYINPUT114), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n762_), .A2(new_n772_), .A3(new_n481_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n520_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n758_), .A2(new_n760_), .A3(new_n749_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n753_), .A2(new_n754_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n774_), .B(new_n481_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT113), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n773_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n742_), .A2(new_n744_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n768_), .A2(new_n769_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n771_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n778_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(new_n780_), .A3(new_n770_), .A4(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n561_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n764_), .A2(KEYINPUT57), .A3(new_n582_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n767_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n576_), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n671_), .B(new_n576_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n487_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(new_n487_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n789_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n392_), .A2(new_n386_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n796_), .A2(new_n258_), .A3(new_n380_), .A4(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n671_), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(KEYINPUT59), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n531_), .A2(new_n247_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(G1340gat));
  NAND3_X1  g604(.A1(new_n801_), .A2(new_n488_), .A3(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n249_), .B1(new_n487_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n799_), .B(new_n808_), .C1(KEYINPUT60), .C2(new_n249_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT116), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(new_n812_), .A3(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1341gat));
  XNOR2_X1  g613(.A(KEYINPUT118), .B(G127gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n803_), .A2(new_n583_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G127gat), .B1(new_n799_), .B2(new_n583_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n818_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n816_), .A2(new_n819_), .A3(new_n820_), .ZN(G1342gat));
  AOI21_X1  g620(.A(G134gat), .B1(new_n799_), .B2(new_n556_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n561_), .A2(G134gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n803_), .B2(new_n823_), .ZN(G1343gat));
  INV_X1    g623(.A(new_n387_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n764_), .B2(new_n582_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n766_), .B(new_n556_), .C1(new_n748_), .C2(new_n763_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n583_), .B1(new_n828_), .B2(new_n786_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n825_), .B(new_n797_), .C1(new_n829_), .C2(new_n794_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n796_), .A2(new_n832_), .A3(new_n825_), .A4(new_n797_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n671_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n488_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n834_), .B2(new_n583_), .ZN(new_n840_));
  AOI211_X1 g639(.A(KEYINPUT120), .B(new_n576_), .C1(new_n831_), .C2(new_n833_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT61), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n387_), .B1(new_n789_), .B2(new_n795_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n832_), .B1(new_n843_), .B2(new_n797_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n794_), .B1(new_n788_), .B2(new_n576_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n797_), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n845_), .A2(KEYINPUT119), .A3(new_n387_), .A4(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n583_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT120), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n834_), .A2(new_n839_), .A3(new_n583_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n842_), .A2(new_n852_), .A3(G155gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(G155gat), .B1(new_n842_), .B2(new_n852_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1346gat));
  AOI21_X1  g654(.A(G162gat), .B1(new_n834_), .B2(new_n556_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n560_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(G162gat), .B2(new_n857_), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n845_), .A2(new_n379_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n257_), .A2(new_n345_), .A3(new_n589_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n671_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G169gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT121), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(new_n864_), .A3(G169gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n865_), .A3(KEYINPUT62), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(KEYINPUT121), .A3(new_n867_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n861_), .A2(new_n307_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT122), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n866_), .A2(new_n868_), .A3(new_n872_), .A4(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1348gat));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n859_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT123), .B1(new_n845_), .B2(new_n379_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n876_), .A2(new_n860_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n488_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G176gat), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n859_), .A2(new_n397_), .A3(new_n488_), .A4(new_n860_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT124), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n884_), .A3(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1349gat));
  AOI21_X1  g685(.A(G183gat), .B1(new_n878_), .B2(new_n583_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n859_), .A2(new_n860_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n888_), .A2(new_n213_), .A3(new_n576_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1350gat));
  OAI21_X1  g689(.A(G190gat), .B1(new_n888_), .B2(new_n560_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n556_), .A2(new_n303_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n888_), .B2(new_n892_), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n345_), .A2(new_n589_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n843_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n671_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g697(.A1(new_n895_), .A2(new_n487_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT125), .B(G204gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1353gat));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n583_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  AND2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n902_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n902_), .B2(new_n903_), .ZN(G1354gat));
  NOR2_X1   g705(.A1(new_n895_), .A2(new_n582_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT126), .ZN(new_n908_));
  INV_X1    g707(.A(G218gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n561_), .A2(G218gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT127), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n908_), .A2(new_n909_), .B1(new_n896_), .B2(new_n911_), .ZN(G1355gat));
endmodule


