//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G232gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G29gat), .B(G36gat), .Z(new_n207_));
  XOR2_X1   g006(.A(G43gat), .B(G50gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT15), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT65), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT7), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n220_), .A2(new_n211_), .A3(new_n212_), .A4(KEYINPUT65), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  OAI22_X1  g028(.A1(new_n223_), .A2(new_n224_), .B1(KEYINPUT9), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G85gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n229_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT64), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n242_), .A2(new_n212_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n237_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n222_), .A2(KEYINPUT66), .A3(KEYINPUT8), .A4(new_n225_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n228_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n210_), .A2(new_n246_), .ZN(new_n247_));
  AOI211_X1 g046(.A(new_n203_), .B(new_n206_), .C1(new_n247_), .C2(KEYINPUT69), .ZN(new_n248_));
  INV_X1    g047(.A(new_n209_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n210_), .B2(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n206_), .A2(new_n203_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n254_), .B2(new_n248_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT70), .ZN(new_n256_));
  XOR2_X1   g055(.A(G190gat), .B(G218gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G134gat), .B(G162gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT36), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n255_), .A2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(KEYINPUT36), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n256_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n256_), .B1(new_n263_), .B2(new_n262_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n202_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n263_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n256_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n256_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT37), .A3(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274_));
  INV_X1    g073(.A(G1gat), .ZN(new_n275_));
  INV_X1    g074(.A(G8gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G8gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G57gat), .B(G64gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G71gat), .B(G78gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT11), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n286_));
  INV_X1    g085(.A(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n283_), .A2(KEYINPUT11), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n285_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n282_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G127gat), .B(G155gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT16), .ZN(new_n293_));
  XOR2_X1   g092(.A(G183gat), .B(G211gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT17), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n296_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n291_), .A2(new_n298_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT71), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(KEYINPUT71), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT72), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n306_), .B(new_n300_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n290_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT12), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n239_), .A2(new_n243_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n313_), .A2(new_n237_), .B1(new_n227_), .B2(new_n226_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n290_), .B1(new_n314_), .B2(new_n245_), .ZN(new_n315_));
  AND4_X1   g114(.A1(new_n245_), .A2(new_n228_), .A3(new_n244_), .A4(new_n290_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n312_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G230gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n246_), .A2(new_n310_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n311_), .ZN(new_n321_));
  AOI211_X1 g120(.A(KEYINPUT67), .B(KEYINPUT12), .C1(new_n246_), .C2(new_n310_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n317_), .B(new_n318_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n315_), .A2(new_n316_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n323_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT5), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  XNOR2_X1  g128(.A(new_n325_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT13), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n273_), .A2(new_n309_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT73), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT89), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT3), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT2), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(KEYINPUT79), .A3(new_n347_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n343_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n340_), .B1(KEYINPUT1), .B2(new_n342_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(KEYINPUT1), .B2(new_n342_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n344_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n346_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G127gat), .B(G134gat), .Z(new_n359_));
  XOR2_X1   g158(.A(G113gat), .B(G120gat), .Z(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(new_n361_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n339_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n369_), .A3(KEYINPUT4), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT90), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n369_), .B2(KEYINPUT4), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n352_), .A2(new_n357_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(KEYINPUT90), .A3(new_n375_), .A4(new_n368_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n370_), .B1(new_n377_), .B2(new_n339_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G57gat), .B(G85gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  AOI211_X1 g184(.A(new_n383_), .B(new_n370_), .C1(new_n377_), .C2(new_n339_), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT96), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT96), .B1(new_n385_), .B2(new_n386_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(G183gat), .A3(G190gat), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(KEYINPUT77), .ZN(new_n393_));
  INV_X1    g192(.A(G183gat), .ZN(new_n394_));
  INV_X1    g193(.A(G190gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT23), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n392_), .A3(KEYINPUT77), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G169gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G169gat), .A2(G176gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n407_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n396_), .A2(new_n392_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(KEYINPUT75), .A2(G183gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT25), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n395_), .A2(KEYINPUT26), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(KEYINPUT76), .A3(G190gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT76), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n413_), .A2(new_n414_), .A3(new_n416_), .A4(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n401_), .A2(new_n403_), .B1(new_n411_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n421_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(new_n368_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427_));
  INV_X1    g226(.A(G15gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT30), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT31), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n426_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n390_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G8gat), .B(G36gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n404_), .B(KEYINPUT85), .Z(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT22), .B(G169gat), .Z(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(G176gat), .ZN(new_n444_));
  AOI211_X1 g243(.A(new_n442_), .B(new_n444_), .C1(new_n410_), .C2(new_n400_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n398_), .A2(new_n409_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT84), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n398_), .A2(new_n448_), .A3(new_n409_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT25), .B(G183gat), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n414_), .A2(new_n417_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n408_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n445_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G211gat), .B(G218gat), .Z(new_n459_));
  INV_X1    g258(.A(KEYINPUT21), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G197gat), .B(G204gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n459_), .A3(KEYINPUT21), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n441_), .B1(new_n458_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT86), .B1(new_n421_), .B2(new_n466_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n463_), .A2(new_n465_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n401_), .A2(new_n403_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n411_), .A2(new_n420_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n472_), .B(new_n473_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n471_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n467_), .A2(new_n477_), .A3(KEYINPUT87), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n441_), .B1(new_n421_), .B2(new_n466_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n458_), .B2(new_n466_), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n470_), .B(KEYINPUT83), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT87), .B1(new_n467_), .B2(new_n477_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n440_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n467_), .A2(new_n477_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n439_), .A3(new_n482_), .A4(new_n478_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n490_), .A2(KEYINPUT27), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n480_), .A2(new_n481_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n458_), .A2(new_n466_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT93), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n456_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n496_), .A2(new_n473_), .A3(new_n445_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n497_), .B2(new_n441_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n471_), .A2(new_n476_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n492_), .B1(new_n500_), .B2(new_n470_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT27), .B(new_n489_), .C1(new_n501_), .C2(new_n439_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n491_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n358_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT80), .B(KEYINPUT28), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G22gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n473_), .A2(KEYINPUT81), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n510_), .A2(G228gat), .A3(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n473_), .B1(new_n358_), .B2(new_n504_), .ZN(new_n513_));
  INV_X1    g312(.A(G78gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(G106gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n513_), .B(G78gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n212_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n512_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n516_), .A2(new_n518_), .A3(new_n512_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n509_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n509_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n519_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n434_), .A2(new_n503_), .A3(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(new_n525_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n385_), .A2(KEYINPUT33), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n385_), .A2(KEYINPUT33), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n365_), .A2(new_n339_), .A3(new_n369_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n384_), .B(new_n531_), .C1(new_n377_), .C2(new_n339_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n490_), .A2(new_n529_), .A3(new_n530_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n439_), .A2(KEYINPUT32), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT92), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n488_), .A2(new_n482_), .A3(new_n478_), .A4(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n470_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n499_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n493_), .A2(KEYINPUT20), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n495_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n543_), .B2(new_n494_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n538_), .B(new_n539_), .C1(new_n544_), .C2(new_n492_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT94), .B1(new_n501_), .B2(new_n534_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n537_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n533_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT95), .B(new_n537_), .C1(new_n546_), .C2(new_n545_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n528_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n526_), .A2(new_n390_), .A3(new_n491_), .A4(new_n502_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n527_), .B1(new_n553_), .B2(new_n432_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n280_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT74), .B1(new_n555_), .B2(new_n209_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n209_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G229gat), .A3(G233gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n210_), .A2(new_n280_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n560_), .B(new_n561_), .C1(new_n249_), .C2(new_n280_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G169gat), .B(G197gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n563_), .B(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n337_), .A2(new_n554_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT38), .ZN(new_n570_));
  AOI21_X1  g369(.A(G1gat), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n389_), .A3(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n569_), .A2(new_n570_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n269_), .A2(new_n270_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n554_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n334_), .A2(new_n567_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n309_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT98), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n389_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n581_), .A2(KEYINPUT99), .A3(G1gat), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT99), .B1(new_n581_), .B2(G1gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n574_), .B1(new_n582_), .B2(new_n583_), .ZN(G1324gat));
  NAND3_X1  g383(.A1(new_n568_), .A2(new_n276_), .A3(new_n503_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n576_), .A2(new_n503_), .A3(new_n579_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  AND4_X1   g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .A4(G8gat), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n276_), .B1(KEYINPUT100), .B2(KEYINPUT39), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n587_), .A2(new_n590_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n585_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(G1325gat));
  NAND3_X1  g393(.A1(new_n568_), .A2(new_n428_), .A3(new_n433_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n580_), .A2(new_n433_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G15gat), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT41), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT41), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n596_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n597_), .A2(new_n600_), .A3(new_n601_), .A4(new_n602_), .ZN(G1326gat));
  INV_X1    g402(.A(G22gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n568_), .A2(new_n604_), .A3(new_n526_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n580_), .A2(new_n526_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G22gat), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT42), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT42), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(G1327gat));
  AOI21_X1  g409(.A(new_n433_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n272_), .B1(new_n611_), .B2(new_n527_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT43), .B(new_n272_), .C1(new_n611_), .C2(new_n527_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n308_), .A3(new_n577_), .A4(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n309_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(KEYINPUT44), .A3(new_n577_), .A4(new_n615_), .ZN(new_n620_));
  AND4_X1   g419(.A1(G29gat), .A2(new_n618_), .A3(new_n389_), .A4(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n554_), .A2(new_n567_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n575_), .A2(new_n308_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT103), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n334_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n389_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n621_), .A2(new_n628_), .ZN(G1328gat));
  NAND3_X1  g428(.A1(new_n618_), .A2(new_n503_), .A3(new_n620_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G36gat), .ZN(new_n631_));
  INV_X1    g430(.A(G36gat), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n622_), .A2(new_n632_), .A3(new_n503_), .A4(new_n625_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT45), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n631_), .A2(KEYINPUT46), .A3(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1329gat));
  NOR2_X1   g438(.A1(new_n432_), .A2(new_n423_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n618_), .A2(new_n620_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n618_), .A2(KEYINPUT104), .A3(new_n620_), .A4(new_n640_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n423_), .B1(new_n626_), .B2(new_n432_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT47), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT47), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n643_), .A2(new_n648_), .A3(new_n644_), .A4(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(G1330gat));
  NAND3_X1  g449(.A1(new_n618_), .A2(new_n526_), .A3(new_n620_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G50gat), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n528_), .A2(G50gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT105), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n627_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT106), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1331gat));
  NAND3_X1  g459(.A1(new_n305_), .A2(new_n307_), .A3(new_n567_), .ZN(new_n661_));
  NOR4_X1   g460(.A1(new_n554_), .A2(new_n575_), .A3(new_n335_), .A4(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(G57gat), .A3(new_n389_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT108), .Z(new_n664_));
  INV_X1    g463(.A(G57gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n554_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT107), .A3(new_n567_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  INV_X1    g467(.A(new_n567_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n554_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n272_), .A2(new_n308_), .A3(new_n335_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n389_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n664_), .B1(new_n665_), .B2(new_n673_), .ZN(G1332gat));
  NAND2_X1  g473(.A1(new_n662_), .A2(new_n503_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G64gat), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT48), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT48), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n671_), .A2(new_n672_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G64gat), .B1(new_n491_), .B2(new_n502_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT109), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n677_), .A2(new_n678_), .B1(new_n679_), .B2(new_n681_), .ZN(G1333gat));
  OR3_X1    g481(.A1(new_n679_), .A2(G71gat), .A3(new_n432_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n662_), .A2(new_n433_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT49), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G71gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G71gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n683_), .B(KEYINPUT110), .C1(new_n687_), .C2(new_n686_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1334gat));
  NAND2_X1  g491(.A1(new_n662_), .A2(new_n526_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G78gat), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT50), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT50), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n526_), .A2(new_n514_), .ZN(new_n697_));
  OAI22_X1  g496(.A1(new_n695_), .A2(new_n696_), .B1(new_n679_), .B2(new_n697_), .ZN(G1335gat));
  AOI211_X1 g497(.A(new_n335_), .B(new_n624_), .C1(new_n667_), .C2(new_n670_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n231_), .A3(new_n389_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n619_), .A2(new_n615_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n335_), .A2(new_n669_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n389_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n704_), .B2(new_n231_), .ZN(G1336gat));
  AOI21_X1  g504(.A(G92gat), .B1(new_n699_), .B2(new_n503_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n503_), .A2(G92gat), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT111), .Z(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n703_), .B2(new_n708_), .ZN(G1337gat));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(KEYINPUT112), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n432_), .A2(new_n241_), .A3(new_n240_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n699_), .B2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n701_), .A2(new_n433_), .A3(new_n702_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G99gat), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n710_), .A2(KEYINPUT112), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(G1338gat));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n212_), .A3(new_n526_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n619_), .A2(new_n526_), .A3(new_n615_), .A4(new_n702_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(G106gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G106gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n724_), .B(new_n726_), .ZN(G1339gat));
  INV_X1    g526(.A(new_n566_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n558_), .A2(new_n561_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n561_), .B1(new_n555_), .B2(new_n209_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n566_), .B1(new_n560_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT119), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n563_), .A2(new_n728_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n733_), .B2(new_n732_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n325_), .A2(new_n329_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n323_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT116), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n323_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n318_), .A2(new_n739_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n317_), .B(new_n745_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(KEYINPUT117), .A2(G230gat), .A3(G233gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n317_), .B(new_n749_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n738_), .B1(new_n744_), .B2(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n323_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n742_), .B1(new_n323_), .B2(new_n739_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n751_), .B(new_n738_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n329_), .B1(new_n752_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT118), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n755_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n329_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n737_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n272_), .B1(new_n764_), .B2(KEYINPUT58), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT120), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(KEYINPUT58), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n272_), .B(new_n768_), .C1(new_n764_), .C2(KEYINPUT58), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n669_), .A2(new_n736_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT56), .B1(new_n762_), .B2(new_n329_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n329_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n758_), .B(new_n773_), .C1(new_n761_), .C2(new_n755_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n735_), .A2(new_n330_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n575_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT57), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n575_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n309_), .B1(new_n770_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n661_), .A2(KEYINPUT114), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n305_), .A2(new_n307_), .A3(new_n786_), .A4(new_n567_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(new_n334_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n335_), .A2(new_n785_), .A3(KEYINPUT115), .A4(new_n787_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n273_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n783_), .A2(new_n793_), .ZN(new_n794_));
  NOR4_X1   g593(.A1(new_n503_), .A2(new_n526_), .A3(new_n390_), .A4(new_n432_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(G113gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n669_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n795_), .C1(new_n783_), .C2(new_n793_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT121), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT121), .B(new_n795_), .C1(new_n783_), .C2(new_n793_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(KEYINPUT59), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n801_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n567_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n798_), .B1(new_n807_), .B2(new_n797_), .ZN(G1340gat));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n335_), .B2(KEYINPUT60), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n796_), .B(new_n810_), .C1(KEYINPUT60), .C2(new_n809_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n335_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n809_), .ZN(G1341gat));
  INV_X1    g612(.A(G127gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n796_), .A2(new_n814_), .A3(new_n309_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n308_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n814_), .ZN(G1342gat));
  INV_X1    g616(.A(G134gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n796_), .A2(new_n818_), .A3(new_n575_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n273_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n818_), .ZN(G1343gat));
  NOR4_X1   g620(.A1(new_n503_), .A2(new_n528_), .A3(new_n390_), .A4(new_n433_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n794_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n669_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n334_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g626(.A1(new_n794_), .A2(new_n822_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n308_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT61), .B(G155gat), .Z(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  OAI21_X1  g630(.A(G162gat), .B1(new_n828_), .B2(new_n273_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n778_), .A2(G162gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n828_), .B2(new_n833_), .ZN(G1347gat));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n434_), .B1(new_n491_), .B2(new_n502_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(new_n669_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n528_), .B(new_n837_), .C1(new_n783_), .C2(new_n793_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n838_), .A2(new_n443_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT62), .B1(new_n838_), .B2(G169gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n835_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n842_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(new_n839_), .A3(KEYINPUT123), .A4(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1348gat));
  OAI211_X1 g645(.A(new_n528_), .B(new_n836_), .C1(new_n783_), .C2(new_n793_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n335_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(G176gat), .Z(G1349gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n308_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n452_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n394_), .B2(new_n850_), .ZN(G1350gat));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n847_), .A2(new_n273_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(G190gat), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n853_), .B(G190gat), .C1(new_n847_), .C2(new_n273_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n575_), .A2(new_n454_), .ZN(new_n858_));
  OAI22_X1  g657(.A1(new_n855_), .A2(new_n857_), .B1(new_n847_), .B2(new_n858_), .ZN(G1351gat));
  AND4_X1   g658(.A1(new_n390_), .A2(new_n503_), .A3(new_n526_), .A4(new_n432_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n794_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n669_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n334_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g664(.A(new_n308_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT125), .Z(new_n867_));
  NOR3_X1   g666(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n870_), .B(new_n872_), .ZN(G1354gat));
  NAND2_X1  g672(.A1(new_n861_), .A2(new_n575_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT127), .B(G218gat), .Z(new_n875_));
  NOR2_X1   g674(.A1(new_n273_), .A2(new_n875_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n875_), .B1(new_n861_), .B2(new_n876_), .ZN(G1355gat));
endmodule


