//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_;
  INV_X1    g000(.A(KEYINPUT9), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(new_n204_), .ZN(new_n209_));
  NAND4_X1  g008(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT10), .B(G99gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n211_), .B(new_n217_), .C1(G106gat), .C2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n223_), .A2(new_n214_), .A3(new_n215_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  XOR2_X1   g025(.A(G85gat), .B(G92gat), .Z(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n226_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n219_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232_));
  INV_X1    g031(.A(G71gat), .ZN(new_n233_));
  INV_X1    g032(.A(G78gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G71gat), .A2(G78gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT11), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT66), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n239_));
  AND2_X1   g038(.A1(G71gat), .A2(G78gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G71gat), .A2(G78gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G57gat), .ZN(new_n243_));
  INV_X1    g042(.A(G64gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G57gat), .A2(G64gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n240_), .A2(new_n241_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT11), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n238_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n248_), .B1(new_n251_), .B2(new_n238_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n232_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n235_), .A2(new_n236_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n255_), .A2(new_n239_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(new_n249_), .B2(KEYINPUT11), .ZN(new_n257_));
  NOR4_X1   g056(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT66), .A4(new_n239_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n238_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT67), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n231_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT64), .Z(new_n265_));
  NOR3_X1   g064(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n225_), .A2(new_n227_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT8), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n218_), .A2(G106gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(new_n216_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n268_), .A2(new_n228_), .B1(new_n270_), .B2(new_n211_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n259_), .A2(KEYINPUT67), .A3(new_n260_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT67), .B1(new_n259_), .B2(new_n260_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n265_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT69), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n266_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT12), .B1(new_n252_), .B2(new_n253_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n271_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n259_), .A2(new_n260_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n231_), .A2(KEYINPUT68), .A3(new_n281_), .A4(KEYINPUT12), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n254_), .A2(new_n231_), .A3(new_n261_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n280_), .B(new_n282_), .C1(new_n284_), .C2(KEYINPUT12), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT70), .B1(new_n277_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n263_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n274_), .A2(KEYINPUT69), .A3(new_n275_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n272_), .A2(new_n273_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT12), .B1(new_n290_), .B2(new_n231_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n280_), .A2(new_n282_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n286_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n265_), .B1(new_n284_), .B2(new_n262_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G204gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G120gat), .B(G148gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT72), .B(G176gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n297_), .A3(new_n304_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT13), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT13), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G169gat), .B(G197gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G43gat), .B(G50gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT73), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G29gat), .B(G36gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n316_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n323_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G15gat), .B(G22gat), .ZN(new_n328_));
  INV_X1    g127(.A(G1gat), .ZN(new_n329_));
  INV_X1    g128(.A(G8gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT14), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G1gat), .B(G8gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n327_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n324_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n326_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(G229gat), .A3(G233gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n315_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n315_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(KEYINPUT79), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT79), .B1(new_n342_), .B2(new_n343_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT26), .B(G190gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n351_), .A2(G183gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT80), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(KEYINPUT80), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n360_), .A2(KEYINPUT23), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n362_));
  INV_X1    g161(.A(new_n360_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n359_), .A2(new_n364_), .A3(new_n366_), .A4(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G169gat), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n376_), .A2(new_n369_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n360_), .A2(KEYINPUT23), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n363_), .B2(new_n362_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G15gat), .B(G43gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n390_), .B(KEYINPUT86), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n389_), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT85), .Z(new_n393_));
  INV_X1    g192(.A(KEYINPUT31), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n350_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n397_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n349_), .A3(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n365_), .B1(new_n371_), .B2(new_n367_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n356_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n352_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n355_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(new_n379_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n380_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n364_), .A2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n377_), .A2(new_n411_), .A3(KEYINPUT92), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT92), .B1(new_n377_), .B2(new_n411_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(G211gat), .A2(G218gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G211gat), .A2(G218gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT21), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G197gat), .B(G204gat), .ZN(new_n420_));
  AOI211_X1 g219(.A(KEYINPUT90), .B(new_n418_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n419_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n403_), .B1(new_n415_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n414_), .A2(KEYINPUT93), .A3(new_n423_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n423_), .A2(new_n382_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n425_), .A2(KEYINPUT20), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT19), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n423_), .B2(new_n382_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n430_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n433_), .B(new_n434_), .C1(new_n423_), .C2(new_n414_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n437_));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  NOR2_X1   g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT3), .ZN(new_n448_));
  INV_X1    g247(.A(G141gat), .ZN(new_n449_));
  INV_X1    g248(.A(G148gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n451_), .B(new_n452_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n454_), .A2(new_n453_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n446_), .B(new_n447_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n446_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G141gat), .A2(G148gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n449_), .A2(new_n450_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(new_n349_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n457_), .A2(new_n349_), .A3(new_n463_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n467_), .A2(KEYINPUT95), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(KEYINPUT95), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n468_), .A2(G225gat), .A3(G233gat), .A4(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G29gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(new_n203_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT0), .B(G57gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n464_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n467_), .B2(KEYINPUT4), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n475_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT33), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n445_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n482_), .A2(new_n475_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n377_), .A2(new_n411_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n424_), .A2(new_n409_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n433_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n430_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(KEYINPUT32), .A3(new_n443_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n487_), .B(new_n493_), .C1(new_n495_), .C2(new_n436_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n485_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n423_), .B1(new_n498_), .B2(new_n464_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G78gat), .B(G106gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G228gat), .A2(G233gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n423_), .B2(KEYINPUT91), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n501_), .B(new_n503_), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n464_), .A2(new_n498_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT89), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G22gat), .B(G50gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n511_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n505_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n497_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n487_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT27), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n520_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n492_), .A2(new_n441_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(KEYINPUT27), .C1(new_n441_), .C2(new_n436_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n402_), .B1(new_n518_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n517_), .ZN(new_n528_));
  NOR4_X1   g327(.A1(new_n401_), .A2(new_n487_), .A3(new_n528_), .A4(new_n524_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n346_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n312_), .B1(new_n530_), .B2(KEYINPUT96), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n327_), .A2(new_n336_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n231_), .A3(new_n325_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n327_), .A2(new_n271_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT34), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n533_), .B(new_n534_), .C1(KEYINPUT35), .C2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  AND3_X1   g342(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n540_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G183gat), .B(G211gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(G127gat), .B(G155gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT78), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(KEYINPUT17), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n281_), .B(new_n334_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT76), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n562_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n557_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT67), .B1(new_n566_), .B2(new_n559_), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n560_), .B(new_n561_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n558_), .ZN(new_n569_));
  OR3_X1    g368(.A1(new_n565_), .A2(new_n569_), .A3(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT75), .B(new_n572_), .C1(new_n544_), .C2(new_n546_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n552_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n526_), .A2(new_n518_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n402_), .A2(new_n517_), .A3(new_n525_), .ZN(new_n577_));
  OAI22_X1  g376(.A1(new_n576_), .A2(new_n402_), .B1(new_n577_), .B2(new_n487_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n346_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n531_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n583_), .A2(new_n329_), .A3(new_n487_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT38), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n586_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n527_), .A2(new_n529_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT98), .B1(new_n589_), .B2(new_n547_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n591_));
  INV_X1    g390(.A(new_n547_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n578_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n344_), .A2(new_n345_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n312_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n593_), .A3(new_n571_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n487_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n587_), .A2(new_n588_), .A3(new_n600_), .A4(new_n601_), .ZN(G1324gat));
  OAI21_X1  g401(.A(G8gat), .B1(new_n596_), .B2(new_n525_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n605_), .B(G8gat), .C1(new_n596_), .C2(new_n525_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n583_), .A2(new_n330_), .A3(new_n524_), .A4(new_n584_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(G1325gat));
  NOR2_X1   g410(.A1(new_n401_), .A2(G15gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n583_), .A2(new_n584_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G15gat), .B1(new_n596_), .B2(new_n401_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n613_), .B1(new_n617_), .B2(new_n618_), .ZN(G1326gat));
  NOR2_X1   g418(.A1(new_n517_), .A2(G22gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n583_), .A2(new_n584_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G22gat), .B1(new_n596_), .B2(new_n517_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT42), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n622_), .A2(KEYINPUT42), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(G1327gat));
  INV_X1    g425(.A(G29gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n552_), .A2(new_n573_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT43), .B1(new_n589_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n578_), .A2(new_n631_), .A3(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n571_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n595_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n571_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(KEYINPUT44), .A3(new_n595_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n487_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n627_), .B1(new_n640_), .B2(KEYINPUT102), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(KEYINPUT102), .B2(new_n640_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n592_), .A2(new_n571_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n531_), .A2(new_n580_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT103), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n531_), .A2(new_n646_), .A3(new_n580_), .A4(new_n643_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n645_), .A2(new_n647_), .A3(new_n627_), .A4(new_n487_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n642_), .A2(new_n648_), .ZN(G1328gat));
  OR2_X1    g448(.A1(new_n525_), .A2(KEYINPUT104), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n525_), .A2(KEYINPUT104), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(G36gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n645_), .A2(new_n647_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT45), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n645_), .A2(new_n647_), .A3(new_n656_), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n637_), .A2(new_n524_), .A3(new_n639_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n660_), .A3(KEYINPUT46), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1329gat));
  NAND4_X1  g464(.A1(new_n637_), .A2(new_n639_), .A3(G43gat), .A4(new_n402_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n645_), .A2(new_n402_), .A3(new_n647_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(G43gat), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g468(.A(G50gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n637_), .A2(new_n528_), .A3(new_n639_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(KEYINPUT105), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(KEYINPUT105), .B2(new_n671_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n645_), .A2(new_n647_), .A3(new_n670_), .A4(new_n528_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1331gat));
  NOR2_X1   g474(.A1(new_n311_), .A2(new_n346_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n578_), .A2(new_n575_), .A3(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT106), .Z(new_n678_));
  AOI21_X1  g477(.A(G57gat), .B1(new_n678_), .B2(new_n487_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n590_), .A2(new_n571_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(new_n593_), .A3(new_n676_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n243_), .A3(new_n597_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1332gat));
  INV_X1    g482(.A(new_n652_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n678_), .A2(new_n244_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G64gat), .B1(new_n681_), .B2(new_n652_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n686_), .A2(KEYINPUT48), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1333gat));
  NAND3_X1  g489(.A1(new_n678_), .A2(new_n233_), .A3(new_n402_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n680_), .A2(new_n402_), .A3(new_n593_), .A4(new_n676_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT49), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(G71gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n692_), .B2(G71gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n691_), .B(KEYINPUT107), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  NAND3_X1  g500(.A1(new_n678_), .A2(new_n234_), .A3(new_n528_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G78gat), .B1(new_n681_), .B2(new_n517_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT50), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n703_), .A2(KEYINPUT50), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1335gat));
  NAND3_X1  g506(.A1(new_n578_), .A2(new_n643_), .A3(new_n676_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n709_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n597_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(KEYINPUT109), .A3(G85gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(KEYINPUT109), .B1(new_n712_), .B2(G85gat), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n638_), .A2(G85gat), .A3(new_n487_), .A4(new_n676_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n713_), .A2(KEYINPUT110), .A3(new_n714_), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1336gat));
  NAND2_X1  g519(.A1(new_n710_), .A2(new_n711_), .ZN(new_n721_));
  AOI21_X1  g520(.A(G92gat), .B1(new_n721_), .B2(new_n524_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT111), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(KEYINPUT111), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n638_), .A2(new_n676_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n725_), .A2(new_n204_), .A3(new_n652_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(G1337gat));
  OAI21_X1  g526(.A(G99gat), .B1(new_n725_), .B2(new_n401_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n401_), .A2(new_n218_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n721_), .A2(KEYINPUT112), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT112), .B1(new_n721_), .B2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n721_), .A2(new_n222_), .A3(new_n528_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n638_), .A2(new_n528_), .A3(new_n676_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G106gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G106gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g539(.A1(new_n577_), .A2(new_n597_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n337_), .A2(new_n338_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n315_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n335_), .B1(G229gat), .B2(G233gat), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n341_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n308_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n289_), .A2(new_n293_), .A3(KEYINPUT55), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n289_), .A2(new_n293_), .A3(new_n753_), .A4(KEYINPUT55), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n293_), .A2(new_n274_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n265_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT55), .B1(new_n286_), .B2(new_n295_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n305_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n289_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n294_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n751_), .A2(KEYINPUT114), .B1(new_n755_), .B2(new_n265_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n754_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n305_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT115), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT56), .B(new_n305_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n307_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n594_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n750_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n743_), .B1(new_n776_), .B2(new_n547_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n346_), .A2(new_n307_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n772_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n762_), .B2(new_n761_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n778_), .B1(new_n780_), .B2(new_n771_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT57), .B(new_n592_), .C1(new_n781_), .C2(new_n750_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n761_), .A2(new_n784_), .A3(new_n772_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n307_), .A2(new_n748_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n761_), .B2(new_n784_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n770_), .B2(KEYINPUT116), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n761_), .A2(new_n784_), .A3(new_n772_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT58), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n628_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n777_), .A2(new_n782_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n634_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n574_), .A2(new_n346_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n311_), .ZN(new_n797_));
  OR2_X1    g596(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n798_));
  NAND2_X1  g597(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n796_), .A2(KEYINPUT113), .A3(KEYINPUT54), .A4(new_n311_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n742_), .B1(new_n795_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G113gat), .B1(new_n804_), .B2(new_n346_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n741_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n772_), .B1(new_n770_), .B2(KEYINPUT115), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n761_), .A2(new_n762_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n775_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n547_), .B1(new_n810_), .B2(new_n749_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n793_), .B(KEYINPUT118), .C1(new_n811_), .C2(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n782_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT118), .B1(new_n777_), .B2(new_n793_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n634_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n807_), .B1(new_n815_), .B2(new_n803_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT117), .B1(new_n804_), .B2(new_n806_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n802_), .B1(new_n794_), .B2(new_n634_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n818_), .B(KEYINPUT59), .C1(new_n819_), .C2(new_n742_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n346_), .A2(G113gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n805_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT119), .B(G120gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n821_), .B2(new_n312_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n311_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n804_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n826_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n824_), .B1(new_n827_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n816_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n592_), .B1(new_n781_), .B2(new_n750_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n790_), .A2(new_n791_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n629_), .B1(new_n835_), .B2(new_n783_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n834_), .A2(new_n743_), .B1(new_n792_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n571_), .B1(new_n837_), .B2(new_n782_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n741_), .B1(new_n838_), .B2(new_n802_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n818_), .B1(new_n839_), .B2(KEYINPUT59), .ZN(new_n840_));
  INV_X1    g639(.A(new_n820_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n833_), .B(new_n312_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n825_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n829_), .B(KEYINPUT120), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(KEYINPUT121), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n832_), .A2(new_n845_), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n804_), .B2(new_n571_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n571_), .A2(G127gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n821_), .B2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n804_), .B2(new_n547_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n628_), .A2(G134gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n821_), .B2(new_n851_), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n819_), .A2(new_n402_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n684_), .A2(new_n597_), .A3(new_n517_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n594_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n449_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n311_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n450_), .ZN(G1345gat));
  INV_X1    g658(.A(new_n855_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n571_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT122), .B1(new_n855_), .B2(new_n634_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n864_), .B(new_n866_), .ZN(G1346gat));
  AND3_X1   g666(.A1(new_n860_), .A2(G162gat), .A3(new_n628_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G162gat), .B1(new_n860_), .B2(new_n547_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1347gat));
  INV_X1    g669(.A(G169gat), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n652_), .A2(new_n487_), .A3(new_n528_), .A4(new_n401_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n815_), .B2(new_n803_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n874_), .B2(new_n346_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n594_), .B(new_n873_), .C1(new_n815_), .C2(new_n803_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n881_), .B(new_n876_), .C1(new_n882_), .C2(new_n871_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT125), .B1(new_n875_), .B2(new_n877_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n875_), .A2(KEYINPUT124), .A3(new_n877_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n880_), .A2(new_n883_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n374_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1348gat));
  INV_X1    g687(.A(new_n819_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n889_), .A2(G176gat), .A3(new_n312_), .A4(new_n872_), .ZN(new_n890_));
  AOI211_X1 g689(.A(KEYINPUT126), .B(G176gat), .C1(new_n874_), .C2(new_n312_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n815_), .A2(new_n803_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n312_), .A3(new_n872_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n894_), .B2(new_n375_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n890_), .B1(new_n891_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT127), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n898_), .B(new_n890_), .C1(new_n891_), .C2(new_n895_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n873_), .A2(new_n634_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G183gat), .B1(new_n889_), .B2(new_n901_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n571_), .A2(new_n406_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n874_), .B2(new_n903_), .ZN(G1350gat));
  INV_X1    g703(.A(new_n874_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G190gat), .B1(new_n905_), .B2(new_n629_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n874_), .A2(new_n547_), .A3(new_n355_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1351gat));
  AND3_X1   g707(.A1(new_n853_), .A2(new_n519_), .A3(new_n684_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n346_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n312_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n571_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AND2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  AOI21_X1  g717(.A(G218gat), .B1(new_n909_), .B2(new_n547_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n628_), .A2(G218gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n909_), .B2(new_n920_), .ZN(G1355gat));
endmodule


