//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n974_, new_n975_, new_n977_, new_n978_,
    new_n979_, new_n981_, new_n982_, new_n983_, new_n984_, new_n986_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n995_, new_n996_, new_n997_, new_n998_;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT75), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(G29gat), .B(G36gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G15gat), .B(G22gat), .ZN(new_n211_));
  INV_X1    g010(.A(G1gat), .ZN(new_n212_));
  INV_X1    g011(.A(G8gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G1gat), .B(G8gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n218_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT74), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n210_), .A2(KEYINPUT74), .A3(new_n218_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n222_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n210_), .B(KEYINPUT15), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(new_n217_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n205_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n205_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT23), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246_));
  INV_X1    g045(.A(G169gat), .ZN(new_n247_));
  INV_X1    g046(.A(G176gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n245_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G183gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT76), .B1(new_n252_), .B2(KEYINPUT25), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(G183gat), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(KEYINPUT25), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n257_), .A2(KEYINPUT77), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n253_), .A2(new_n256_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n251_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n239_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT79), .B1(new_n247_), .B2(KEYINPUT22), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(G169gat), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n267_), .A2(new_n270_), .A3(new_n248_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n247_), .A2(KEYINPUT78), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n247_), .A2(KEYINPUT78), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT22), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n266_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n242_), .A2(new_n244_), .A3(KEYINPUT80), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT80), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n241_), .A2(new_n277_), .A3(KEYINPUT23), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n278_), .C1(G183gat), .C2(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n265_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT30), .B1(new_n265_), .B2(new_n280_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n236_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND4_X1   g084(.A1(new_n258_), .A2(new_n259_), .A3(new_n256_), .A4(new_n253_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n250_), .B1(new_n286_), .B2(KEYINPUT77), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n287_), .A2(new_n264_), .B1(new_n279_), .B2(new_n275_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT30), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n281_), .A2(new_n282_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n236_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G227gat), .A2(G233gat), .ZN(new_n293_));
  INV_X1    g092(.A(G15gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G43gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT83), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n285_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n302_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT82), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT31), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n298_), .A2(new_n299_), .B1(new_n300_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n285_), .A2(new_n292_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n297_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n309_), .A2(new_n300_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n285_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(KEYINPUT83), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT84), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n310_), .A2(new_n316_), .A3(new_n320_), .A4(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328_));
  INV_X1    g127(.A(G141gat), .ZN(new_n329_));
  INV_X1    g128(.A(G148gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  NOR3_X1   g131(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n331_), .B(new_n332_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n333_), .A2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n327_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338_));
  XOR2_X1   g137(.A(G141gat), .B(G148gat), .Z(new_n339_));
  NAND3_X1  g138(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n340_), .C1(KEYINPUT1), .C2(new_n326_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n308_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n337_), .A2(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT86), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n308_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n303_), .A2(new_n305_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n325_), .B(new_n346_), .C1(new_n353_), .C2(new_n345_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n350_), .A2(new_n352_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n324_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n344_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n348_), .A2(new_n349_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G22gat), .B(G50gat), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n365_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT28), .B1(new_n344_), .B2(KEYINPUT29), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G197gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT88), .B1(new_n377_), .B2(G204gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(G204gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n377_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT21), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n377_), .B2(G204gat), .ZN(new_n384_));
  INV_X1    g183(.A(G204gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT21), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n384_), .A2(new_n386_), .A3(new_n387_), .A4(new_n379_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G211gat), .B(G218gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n382_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n387_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(new_n379_), .A3(new_n386_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT87), .B1(new_n344_), .B2(KEYINPUT29), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n348_), .A2(KEYINPUT29), .A3(new_n349_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n397_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n347_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n395_), .B1(new_n406_), .B2(new_n394_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n402_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n344_), .A2(KEYINPUT87), .A3(KEYINPUT29), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n399_), .A2(new_n400_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n396_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n403_), .B1(new_n412_), .B2(new_n407_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n376_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n371_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n375_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n409_), .A2(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n364_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n245_), .B1(G183gat), .B2(G190gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT22), .B(G169gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n266_), .B1(new_n422_), .B2(new_n248_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT26), .B(G190gat), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n255_), .A2(G183gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n259_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n240_), .B(new_n249_), .C1(new_n425_), .C2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n276_), .A2(new_n278_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n424_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n420_), .B1(new_n394_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT19), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n388_), .A2(new_n389_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n435_), .A2(new_n382_), .B1(new_n392_), .B2(new_n391_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n265_), .A3(new_n280_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n434_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n239_), .A2(KEYINPUT24), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n249_), .B1(new_n440_), .B2(new_n237_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n427_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n258_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n429_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n443_), .A2(new_n444_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n420_), .B1(new_n445_), .B2(new_n436_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT91), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n281_), .A2(new_n447_), .A3(new_n394_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n281_), .B2(new_n394_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n446_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n439_), .B1(new_n450_), .B2(new_n433_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G8gat), .B(G36gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n419_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n446_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT91), .B1(new_n288_), .B2(new_n436_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n281_), .A2(new_n447_), .A3(new_n394_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n438_), .B1(new_n460_), .B2(new_n434_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n455_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(KEYINPUT95), .A3(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n433_), .A2(new_n420_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n445_), .A2(new_n436_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(KEYINPUT92), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n445_), .A2(new_n436_), .A3(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n467_), .B(new_n469_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT93), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n431_), .A2(new_n437_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n433_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n458_), .A2(new_n459_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT92), .B1(new_n394_), .B2(new_n430_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n475_), .A2(new_n469_), .A3(new_n464_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(new_n473_), .A3(new_n478_), .A4(new_n455_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n456_), .A2(new_n463_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT27), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n473_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n477_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n462_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT27), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n479_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n418_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n409_), .A2(new_n413_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n376_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n376_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n461_), .A2(KEYINPUT32), .A3(new_n455_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n455_), .A2(KEYINPUT32), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT94), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n471_), .A2(new_n496_), .A3(new_n473_), .A4(new_n478_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n493_), .B(new_n497_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n324_), .B(new_n346_), .C1(new_n353_), .C2(new_n345_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n360_), .B1(new_n355_), .B2(new_n325_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n361_), .A2(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT33), .A4(new_n360_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(new_n484_), .A3(new_n479_), .A4(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n492_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n323_), .B1(new_n487_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n481_), .A2(new_n486_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n414_), .A2(new_n417_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n507_), .A2(new_n322_), .A3(new_n364_), .A4(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n235_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(G85gat), .B(G92gat), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT6), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(G99gat), .A3(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  INV_X1    g320(.A(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n515_), .A2(new_n520_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G85gat), .B(G92gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n517_), .A2(new_n519_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530_));
  INV_X1    g329(.A(G99gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n522_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n528_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT8), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n518_), .B1(G99gat), .B2(G106gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n516_), .A2(KEYINPUT6), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n533_), .B(new_n532_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n528_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n526_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n210_), .A2(new_n542_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n210_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n533_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AOI211_X1 g351(.A(KEYINPUT8), .B(new_n527_), .C1(new_n552_), .C2(new_n520_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n540_), .B1(new_n539_), .B2(new_n528_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT67), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n536_), .A2(new_n556_), .A3(new_n541_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n526_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n547_), .B1(new_n549_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n546_), .A2(new_n543_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n560_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n566_), .B(new_n547_), .C1(new_n549_), .C2(new_n558_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n564_), .B(KEYINPUT36), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n561_), .B2(new_n567_), .ZN(new_n572_));
  OR3_X1    g371(.A1(new_n569_), .A2(KEYINPUT37), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT37), .B1(new_n569_), .B2(new_n572_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT72), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n217_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT73), .ZN(new_n579_));
  INV_X1    g378(.A(G71gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(G78gat), .ZN(new_n581_));
  INV_X1    g380(.A(G78gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(G71gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n585_), .B2(KEYINPUT11), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT65), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n585_), .B2(KEYINPUT11), .ZN(new_n588_));
  INV_X1    g387(.A(G64gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(G57gat), .ZN(new_n590_));
  INV_X1    g389(.A(G57gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(G64gat), .ZN(new_n592_));
  AND4_X1   g391(.A1(new_n587_), .A2(new_n590_), .A3(new_n592_), .A4(KEYINPUT11), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n586_), .B1(new_n588_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n592_), .A3(KEYINPUT11), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT65), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n592_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT11), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n590_), .A2(new_n592_), .A3(new_n587_), .A4(KEYINPUT11), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n596_), .A2(new_n599_), .A3(new_n584_), .A4(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n579_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n604_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n579_), .A2(new_n603_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n609_), .B(new_n605_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n594_), .A2(new_n601_), .A3(KEYINPUT66), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT66), .B1(new_n594_), .B2(new_n601_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n613_), .B1(new_n616_), .B2(new_n578_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n616_), .B2(new_n578_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n575_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT67), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n556_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n525_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n603_), .A2(KEYINPUT12), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n542_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT66), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n602_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n525_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n594_), .A2(new_n601_), .A3(KEYINPUT66), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .A4(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n629_), .A2(new_n634_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n628_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(G120gat), .B(G148gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT5), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n639_), .B(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n647_), .B2(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n621_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n510_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n362_), .A2(new_n363_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n212_), .A3(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT38), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n650_), .A2(new_n235_), .A3(new_n619_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n569_), .A2(KEYINPUT96), .A3(new_n572_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT96), .B1(new_n569_), .B2(new_n572_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n654_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n507_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n504_), .A2(new_n498_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n508_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n322_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n509_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n661_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT97), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n507_), .A2(new_n662_), .B1(new_n664_), .B2(new_n508_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n509_), .B1(new_n671_), .B2(new_n322_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT97), .A3(new_n661_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n658_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n364_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT98), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT98), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n656_), .B1(new_n677_), .B2(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(new_n507_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n659_), .A2(new_n660_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n669_), .B(new_n681_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT97), .B1(new_n672_), .B2(new_n661_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n680_), .B(new_n657_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G8gat), .B1(new_n684_), .B2(KEYINPUT99), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n674_), .B2(new_n680_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT39), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n674_), .A2(new_n686_), .A3(new_n680_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n684_), .A2(KEYINPUT99), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT39), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .A4(G8gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n652_), .A2(G8gat), .A3(new_n507_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT101), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(new_n698_), .A3(new_n695_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n697_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT101), .B(new_n694_), .C1(new_n688_), .C2(new_n692_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n705_), .ZN(G1325gat));
  NAND2_X1  g505(.A1(new_n674_), .A2(new_n322_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(G15gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n707_), .B2(G15gat), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n653_), .A2(new_n294_), .A3(new_n322_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(G1326gat));
  XNOR2_X1  g515(.A(new_n492_), .B(KEYINPUT103), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n652_), .A2(G22gat), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G22gat), .B1(new_n675_), .B2(new_n718_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT42), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT42), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(G1327gat));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  INV_X1    g523(.A(new_n575_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n672_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n672_), .A2(KEYINPUT104), .A3(new_n724_), .A4(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n672_), .A2(new_n725_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT43), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n728_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n650_), .A2(new_n235_), .A3(new_n620_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736_), .B2(new_n364_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n569_), .A2(new_n572_), .ZN(new_n738_));
  AND4_X1   g537(.A1(new_n738_), .A2(new_n510_), .A3(new_n649_), .A4(new_n619_), .ZN(new_n739_));
  INV_X1    g538(.A(G29gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n654_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT105), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1328gat));
  OAI21_X1  g545(.A(G36gat), .B1(new_n736_), .B2(new_n507_), .ZN(new_n747_));
  INV_X1    g546(.A(G36gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n739_), .A2(new_n748_), .A3(new_n680_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT45), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n747_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1329gat));
  XOR2_X1   g553(.A(KEYINPUT107), .B(G43gat), .Z(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n739_), .B2(new_n322_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n734_), .B(KEYINPUT44), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n322_), .A2(G43gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n739_), .B2(new_n717_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n492_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n757_), .B2(new_n762_), .ZN(G1331gat));
  AOI21_X1  g562(.A(new_n234_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(new_n650_), .A3(new_n620_), .A4(new_n575_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT108), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n591_), .A3(new_n654_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n650_), .A2(new_n235_), .A3(new_n620_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n364_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n767_), .A2(new_n771_), .ZN(G1332gat));
  NAND3_X1  g571(.A1(new_n766_), .A2(new_n589_), .A3(new_n680_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G64gat), .B1(new_n770_), .B2(new_n507_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT48), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT48), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n775_), .B2(new_n776_), .ZN(G1333gat));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n580_), .A3(new_n322_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G71gat), .B1(new_n770_), .B2(new_n323_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT49), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT49), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(G1334gat));
  NAND3_X1  g581(.A1(new_n766_), .A2(new_n582_), .A3(new_n717_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G78gat), .B1(new_n770_), .B2(new_n718_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(KEYINPUT50), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(KEYINPUT50), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n785_), .B2(new_n786_), .ZN(G1335gat));
  NOR3_X1   g586(.A1(new_n649_), .A2(new_n234_), .A3(new_n620_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n732_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789_), .B2(new_n364_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n738_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n649_), .A2(new_n791_), .A3(new_n620_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n764_), .A2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n364_), .A2(G85gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(G1336gat));
  INV_X1    g594(.A(G92gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n793_), .B2(new_n507_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT109), .Z(new_n798_));
  NOR3_X1   g597(.A1(new_n789_), .A2(new_n796_), .A3(new_n507_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(G1337gat));
  INV_X1    g599(.A(new_n793_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(new_n322_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT110), .Z(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  OAI21_X1  g603(.A(G99gat), .B1(new_n789_), .B2(new_n323_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n732_), .A2(new_n492_), .A3(new_n788_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n732_), .A2(KEYINPUT112), .A3(new_n492_), .A4(new_n788_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G106gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n809_), .A2(new_n810_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .A4(new_n812_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n793_), .A2(G106gat), .A3(new_n508_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n808_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n808_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n819_), .B(new_n822_), .C1(new_n814_), .C2(new_n817_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1339gat));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n651_), .A2(new_n235_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n651_), .A2(new_n235_), .A3(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n628_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n629_), .B1(new_n558_), .B2(new_n625_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n635_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n616_), .B2(new_n632_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n836_), .A2(new_n637_), .A3(KEYINPUT55), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n833_), .A2(new_n835_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n628_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n837_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n643_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT56), .B(new_n643_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n844_), .A2(KEYINPUT117), .A3(new_n845_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n223_), .B(new_n220_), .C1(new_n549_), .C2(new_n218_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n221_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n205_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n233_), .A2(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n639_), .A2(new_n643_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n849_), .A2(new_n850_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n857_), .A2(new_n858_), .A3(KEYINPUT58), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT58), .B1(new_n857_), .B2(new_n858_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n725_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n234_), .A2(new_n855_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n837_), .A2(new_n841_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT115), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n837_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT56), .B1(new_n868_), .B2(new_n643_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n848_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n854_), .A2(new_n644_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n738_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n862_), .B1(new_n873_), .B2(KEYINPUT57), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n863_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n872_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n791_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(KEYINPUT116), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n874_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n873_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n861_), .A2(new_n880_), .A3(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n831_), .B1(new_n885_), .B2(new_n619_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n323_), .A2(new_n364_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n507_), .A2(new_n508_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n886_), .A2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n825_), .B1(new_n891_), .B2(new_n235_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT120), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n825_), .C1(new_n891_), .C2(new_n235_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT59), .B1(new_n886_), .B2(new_n890_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n890_), .A2(KEYINPUT59), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n873_), .A2(KEYINPUT57), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n850_), .A2(new_n856_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n858_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n857_), .A2(new_n858_), .A3(KEYINPUT58), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n898_), .B1(new_n905_), .B2(new_n725_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n620_), .B1(new_n906_), .B2(new_n884_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n897_), .B1(new_n907_), .B2(new_n831_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n896_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n235_), .A2(new_n825_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n893_), .A2(new_n895_), .B1(new_n909_), .B2(new_n910_), .ZN(G1340gat));
  NAND3_X1  g710(.A1(new_n896_), .A2(new_n650_), .A3(new_n908_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n896_), .A2(KEYINPUT122), .A3(new_n908_), .A4(new_n650_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(G120gat), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n886_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918_));
  AOI21_X1  g717(.A(KEYINPUT121), .B1(new_n918_), .B2(G120gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(G120gat), .B1(new_n650_), .B2(new_n918_), .ZN(new_n920_));
  MUX2_X1   g719(.A(new_n919_), .B(KEYINPUT121), .S(new_n920_), .Z(new_n921_));
  NAND4_X1  g720(.A1(new_n917_), .A2(new_n889_), .A3(new_n887_), .A4(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n922_), .ZN(G1341gat));
  NAND3_X1  g722(.A1(new_n896_), .A2(new_n620_), .A3(new_n908_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G127gat), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n619_), .A2(G127gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n891_), .B2(new_n926_), .ZN(G1342gat));
  NAND3_X1  g726(.A1(new_n896_), .A2(new_n725_), .A3(new_n908_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G134gat), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n661_), .A2(G134gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n891_), .B2(new_n930_), .ZN(G1343gat));
  NOR2_X1   g730(.A1(new_n886_), .A2(new_n322_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n680_), .A2(new_n364_), .A3(new_n508_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n935_), .A2(new_n329_), .A3(new_n234_), .ZN(new_n936_));
  OAI21_X1  g735(.A(G141gat), .B1(new_n934_), .B2(new_n235_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1344gat));
  NAND3_X1  g737(.A1(new_n935_), .A2(new_n330_), .A3(new_n650_), .ZN(new_n939_));
  OAI21_X1  g738(.A(G148gat), .B1(new_n934_), .B2(new_n649_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1345gat));
  XNOR2_X1  g740(.A(KEYINPUT61), .B(G155gat), .ZN(new_n942_));
  OR3_X1    g741(.A1(new_n934_), .A2(new_n619_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n934_), .B2(new_n619_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1346gat));
  OR3_X1    g744(.A1(new_n934_), .A2(G162gat), .A3(new_n661_), .ZN(new_n946_));
  OAI21_X1  g745(.A(G162gat), .B1(new_n934_), .B2(new_n575_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n907_), .A2(new_n831_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n323_), .A2(new_n507_), .A3(new_n654_), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(KEYINPUT123), .Z(new_n951_));
  NOR2_X1   g750(.A1(new_n951_), .A2(new_n717_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT124), .B1(new_n949_), .B2(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n898_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n861_), .A2(new_n955_), .A3(new_n884_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n619_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n831_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n953_), .B1(new_n957_), .B2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n954_), .A2(new_n961_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n962_), .A2(new_n422_), .A3(new_n234_), .ZN(new_n963_));
  AOI211_X1 g762(.A(KEYINPUT62), .B(new_n247_), .C1(new_n959_), .C2(new_n234_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n959_), .A2(new_n234_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n966_), .B2(G169gat), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n963_), .B1(new_n964_), .B2(new_n967_), .ZN(G1348gat));
  INV_X1    g767(.A(new_n951_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n969_), .A2(G176gat), .A3(new_n650_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n886_), .A2(new_n492_), .A3(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n962_), .A2(new_n650_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(new_n248_), .ZN(G1349gat));
  NOR2_X1   g772(.A1(new_n619_), .A2(new_n442_), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n917_), .A2(new_n508_), .A3(new_n620_), .A4(new_n969_), .ZN(new_n975_));
  AOI22_X1  g774(.A1(new_n962_), .A2(new_n974_), .B1(new_n252_), .B2(new_n975_), .ZN(G1350gat));
  NAND3_X1  g775(.A1(new_n962_), .A2(new_n258_), .A3(new_n681_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n575_), .B1(new_n954_), .B2(new_n961_), .ZN(new_n978_));
  INV_X1    g777(.A(G190gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n977_), .B1(new_n978_), .B2(new_n979_), .ZN(G1351gat));
  NOR2_X1   g779(.A1(new_n507_), .A2(new_n418_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n981_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n886_), .A2(new_n322_), .A3(new_n982_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(new_n234_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g784(.A1(new_n983_), .A2(new_n650_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n385_), .A2(KEYINPUT125), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n986_), .B(new_n987_), .ZN(G1353gat));
  AOI21_X1  g787(.A(new_n619_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n989_));
  XOR2_X1   g788(.A(new_n989_), .B(KEYINPUT126), .Z(new_n990_));
  INV_X1    g789(.A(new_n990_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n983_), .A2(new_n991_), .ZN(new_n992_));
  NOR2_X1   g791(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n993_));
  XOR2_X1   g792(.A(new_n992_), .B(new_n993_), .Z(G1354gat));
  AND3_X1   g793(.A1(new_n983_), .A2(G218gat), .A3(new_n725_), .ZN(new_n995_));
  NOR4_X1   g794(.A1(new_n886_), .A2(new_n322_), .A3(new_n661_), .A4(new_n982_), .ZN(new_n996_));
  OR2_X1    g795(.A1(new_n996_), .A2(KEYINPUT127), .ZN(new_n997_));
  AOI21_X1  g796(.A(G218gat), .B1(new_n996_), .B2(KEYINPUT127), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n995_), .B1(new_n997_), .B2(new_n998_), .ZN(G1355gat));
endmodule


