//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n204_), .A2(new_n207_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT65), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n209_), .B2(new_n211_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT65), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n226_));
  AND2_X1   g025(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(new_n226_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  MUX2_X1   g028(.A(new_n226_), .B(new_n228_), .S(new_n229_), .Z(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n217_), .B1(new_n231_), .B2(new_n203_), .ZN(new_n232_));
  AOI211_X1 g031(.A(KEYINPUT8), .B(new_n202_), .C1(new_n230_), .C2(new_n212_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n216_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OR3_X1    g038(.A1(new_n234_), .A2(new_n235_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n238_), .B(KEYINPUT15), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT35), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G232gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT34), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n234_), .A2(new_n241_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n235_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n245_), .A2(new_n242_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G190gat), .B(G218gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G134gat), .B(G162gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(KEYINPUT36), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n240_), .A2(new_n246_), .A3(new_n247_), .A4(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n250_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n253_), .B(KEYINPUT36), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n250_), .B2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT37), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT71), .B(KEYINPUT37), .C1(new_n257_), .C2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n250_), .A2(new_n256_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT72), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n258_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n250_), .A2(KEYINPUT72), .A3(new_n256_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n262_), .A2(new_n263_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G15gat), .B(G22gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(G1gat), .A2(G8gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(KEYINPUT14), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT73), .ZN(new_n274_));
  XOR2_X1   g073(.A(G1gat), .B(G8gat), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n273_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G231gat), .ZN(new_n282_));
  INV_X1    g081(.A(G233gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n276_), .A2(new_n280_), .A3(G231gat), .A4(G233gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G71gat), .B(G78gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(KEYINPUT11), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n290_), .A3(KEYINPUT11), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n288_), .B2(KEYINPUT11), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT67), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n287_), .A4(new_n291_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n298_), .A3(KEYINPUT69), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n298_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n286_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G155gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G183gat), .B(G211gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT17), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n302_), .A2(new_n299_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n284_), .A2(new_n285_), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n303_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n308_), .B(new_n309_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n300_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n286_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n284_), .A2(new_n285_), .A3(new_n316_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n314_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI211_X1 g121(.A(KEYINPUT75), .B(new_n314_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n313_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT76), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT5), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  NAND3_X1  g128(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n311_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n316_), .B2(new_n234_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G230gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT12), .B1(new_n316_), .B2(new_n234_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n316_), .A2(new_n234_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n316_), .A2(new_n234_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n332_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n329_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n334_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n341_), .A2(new_n337_), .A3(new_n332_), .A4(new_n330_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n338_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n333_), .B1(new_n343_), .B2(new_n336_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n329_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT13), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n340_), .A2(KEYINPUT13), .A3(new_n346_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n270_), .A2(new_n325_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G229gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n276_), .A2(new_n280_), .A3(new_n238_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n238_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n354_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n276_), .A2(new_n280_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n241_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n355_), .B(new_n353_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G113gat), .B(G141gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G169gat), .B(G197gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n358_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT77), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n358_), .A2(new_n361_), .A3(new_n367_), .A4(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n358_), .A2(new_n361_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n364_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G169gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT22), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT22), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G169gat), .ZN(new_n377_));
  INV_X1    g176(.A(G176gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT80), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT22), .B(G169gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n378_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(KEYINPUT79), .A2(G183gat), .A3(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT79), .B1(G183gat), .B2(G190gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT23), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT78), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(G169gat), .A3(G176gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n384_), .A2(new_n393_), .A3(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT25), .B(G183gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT26), .B(G190gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n374_), .A2(new_n378_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n395_), .A2(new_n397_), .A3(new_n405_), .A4(KEYINPUT24), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n390_), .A2(KEYINPUT23), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n390_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT23), .B1(new_n410_), .B2(new_n385_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n404_), .B(new_n406_), .C1(new_n408_), .C2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n400_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n413_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(G15gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT30), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n416_), .B(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(KEYINPUT81), .ZN(new_n422_));
  XOR2_X1   g221(.A(G127gat), .B(G134gat), .Z(new_n423_));
  XOR2_X1   g222(.A(G113gat), .B(G120gat), .Z(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT31), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n421_), .A2(KEYINPUT81), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n421_), .A2(KEYINPUT81), .A3(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT19), .ZN(new_n433_));
  INV_X1    g232(.A(G218gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G211gat), .ZN(new_n435_));
  INV_X1    g234(.A(G211gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G218gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT21), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G197gat), .B(G204gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G204gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G197gat), .ZN(new_n443_));
  INV_X1    g242(.A(G197gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G204gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(KEYINPUT21), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n440_), .A2(new_n439_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n441_), .A2(new_n449_), .B1(new_n438_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n400_), .A2(new_n451_), .A3(new_n412_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n389_), .B1(new_n411_), .B2(new_n408_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n398_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n392_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n410_), .A2(new_n385_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(KEYINPUT23), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n394_), .A2(KEYINPUT24), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT90), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT90), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n394_), .A2(new_n461_), .A3(KEYINPUT24), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n405_), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(new_n404_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n441_), .A2(new_n449_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n450_), .A2(new_n438_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n455_), .A2(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT20), .B(new_n452_), .C1(new_n467_), .C2(KEYINPUT91), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n455_), .A2(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n466_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n469_), .A2(KEYINPUT91), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n433_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G8gat), .B(G36gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT18), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G64gat), .B(G92gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT32), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n413_), .A2(new_n470_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n433_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n451_), .A2(new_n455_), .A3(new_n464_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n478_), .A2(KEYINPUT20), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n472_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT92), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n452_), .A2(KEYINPUT20), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n469_), .A2(new_n470_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n467_), .A2(KEYINPUT91), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n484_), .A2(new_n487_), .A3(new_n479_), .A4(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n478_), .A2(KEYINPUT20), .A3(new_n480_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n433_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n477_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n483_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(KEYINPUT92), .A3(new_n493_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G141gat), .A2(G148gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT85), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G141gat), .A2(G148gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT2), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT2), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(G141gat), .A3(G148gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(G141gat), .A2(G148gat), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n503_), .A2(new_n505_), .B1(new_n506_), .B2(KEYINPUT3), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT85), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n497_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n501_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(G155gat), .A2(G162gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G155gat), .A2(G162gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(KEYINPUT86), .A3(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n497_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT1), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(new_n522_), .A3(new_n512_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n524_), .A2(new_n502_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT83), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n521_), .A2(new_n523_), .A3(new_n528_), .A4(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n516_), .A2(new_n517_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n425_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n514_), .A2(new_n515_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n425_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n517_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G225gat), .A2(G233gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G1gat), .B(G29gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G85gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT0), .B(G57gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  AND3_X1   g340(.A1(new_n532_), .A2(KEYINPUT4), .A3(new_n535_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n531_), .A2(new_n543_), .A3(new_n425_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n536_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n537_), .B(new_n541_), .C1(new_n542_), .C2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n532_), .A2(KEYINPUT4), .A3(new_n535_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n545_), .A3(new_n544_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n541_), .B1(new_n550_), .B2(new_n537_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n495_), .B(new_n496_), .C1(new_n548_), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT33), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n472_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n476_), .B1(new_n472_), .B2(new_n481_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n550_), .A2(KEYINPUT33), .A3(new_n537_), .A4(new_n541_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n536_), .A3(new_n544_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n541_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n532_), .A2(new_n535_), .A3(new_n545_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n554_), .A2(new_n557_), .A3(new_n558_), .A4(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G22gat), .B(G50gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G78gat), .B(G106gat), .ZN(new_n565_));
  INV_X1    g364(.A(G228gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT88), .B1(new_n566_), .B2(new_n283_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n565_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n531_), .A2(KEYINPUT29), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n566_), .A2(new_n283_), .A3(KEYINPUT88), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n470_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  AOI211_X1 g373(.A(new_n572_), .B(new_n568_), .C1(new_n531_), .C2(KEYINPUT29), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n564_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT28), .B1(new_n531_), .B2(KEYINPUT29), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT28), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n533_), .A2(new_n578_), .A3(new_n579_), .A4(new_n517_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT89), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT89), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n533_), .B2(new_n517_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n568_), .B1(new_n585_), .B2(new_n572_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n570_), .A2(new_n573_), .A3(new_n569_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n564_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n576_), .A2(new_n582_), .A3(new_n584_), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n582_), .A2(new_n584_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n574_), .A2(new_n575_), .A3(new_n564_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n588_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n552_), .A2(new_n563_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT27), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n472_), .A2(new_n476_), .A3(new_n481_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n489_), .A2(new_n491_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT27), .B(new_n598_), .C1(new_n599_), .C2(new_n476_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n594_), .A2(new_n597_), .A3(new_n590_), .A4(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n548_), .A2(new_n551_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n431_), .B1(new_n595_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n597_), .A2(new_n600_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n594_), .A2(new_n590_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n429_), .A2(new_n430_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n602_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT93), .B(new_n431_), .C1(new_n595_), .C2(new_n603_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n606_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n352_), .A2(new_n373_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(G1gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n602_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT94), .Z(new_n622_));
  INV_X1    g421(.A(new_n268_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n616_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n351_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(KEYINPUT95), .A3(new_n373_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n627_));
  INV_X1    g426(.A(new_n373_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n351_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n324_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n624_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n618_), .B1(new_n633_), .B2(new_n602_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n620_), .B2(new_n619_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n622_), .A2(new_n635_), .ZN(G1324gat));
  XNOR2_X1  g435(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n608_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(G8gat), .ZN(new_n640_));
  INV_X1    g439(.A(G8gat), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT39), .B(new_n641_), .C1(new_n633_), .C2(new_n608_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n617_), .A2(new_n641_), .A3(new_n608_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n637_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n644_), .B(new_n637_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n632_), .B2(new_n431_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT41), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n617_), .A2(new_n418_), .A3(new_n612_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n617_), .A2(new_n653_), .A3(new_n610_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n633_), .A2(new_n610_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(G22gat), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT42), .B(new_n653_), .C1(new_n633_), .C2(new_n610_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT76), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n324_), .B(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n630_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n552_), .A2(new_n563_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n609_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n601_), .A2(new_n602_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT93), .B1(new_n670_), .B2(new_n431_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n615_), .A2(new_n614_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n666_), .B(new_n270_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n666_), .B1(new_n616_), .B2(new_n270_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n665_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n665_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n602_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n662_), .B1(new_n681_), .B2(G29gat), .ZN(new_n682_));
  INV_X1    g481(.A(G29gat), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT98), .B(new_n683_), .C1(new_n680_), .C2(new_n602_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n664_), .A2(new_n623_), .A3(new_n351_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n616_), .A3(new_n373_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT99), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT99), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n602_), .A2(new_n683_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT100), .Z(new_n691_));
  OAI22_X1  g490(.A1(new_n682_), .A2(new_n684_), .B1(new_n689_), .B2(new_n691_), .ZN(G1328gat));
  NOR2_X1   g491(.A1(new_n607_), .A2(G36gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n687_), .A2(new_n688_), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n678_), .A2(new_n608_), .A3(new_n679_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT101), .B1(new_n696_), .B2(G36gat), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT46), .B(new_n695_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n694_), .B(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n696_), .A2(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n699_), .B1(new_n706_), .B2(new_n707_), .ZN(G1329gat));
  NAND4_X1  g507(.A1(new_n678_), .A2(G43gat), .A3(new_n612_), .A4(new_n679_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n689_), .A2(new_n431_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G43gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g511(.A1(new_n689_), .A2(new_n609_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(G50gat), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n610_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n680_), .B2(new_n715_), .ZN(G1331gat));
  AND2_X1   g515(.A1(new_n616_), .A2(new_n628_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n266_), .A2(new_n267_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n250_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n269_), .A3(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n250_), .A2(new_n256_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n258_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT71), .B1(new_n723_), .B2(KEYINPUT37), .ZN(new_n724_));
  INV_X1    g523(.A(new_n263_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n664_), .A3(new_n351_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n717_), .B1(new_n718_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n718_), .B2(new_n727_), .ZN(new_n729_));
  INV_X1    g528(.A(G57gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n602_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n624_), .A2(new_n628_), .A3(new_n664_), .A4(new_n351_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n613_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1332gat));
  OAI21_X1  g533(.A(G64gat), .B1(new_n732_), .B2(new_n607_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT48), .ZN(new_n736_));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n729_), .A2(new_n737_), .A3(new_n608_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1333gat));
  OAI21_X1  g538(.A(G71gat), .B1(new_n732_), .B2(new_n431_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT104), .B(KEYINPUT49), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n729_), .A2(new_n743_), .A3(new_n612_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1334gat));
  OAI21_X1  g544(.A(G78gat), .B1(new_n732_), .B2(new_n609_), .ZN(new_n746_));
  XOR2_X1   g545(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G78gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n729_), .A2(new_n749_), .A3(new_n610_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1335gat));
  OR2_X1    g550(.A1(new_n674_), .A2(new_n675_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n664_), .A2(new_n373_), .A3(new_n625_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT106), .ZN(new_n755_));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n613_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n664_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n717_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(new_n213_), .A3(new_n602_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n756_), .A2(new_n760_), .ZN(G1336gat));
  OAI21_X1  g560(.A(G92gat), .B1(new_n755_), .B2(new_n607_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n214_), .A3(new_n608_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n612_), .A3(new_n205_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n752_), .A2(new_n612_), .A3(new_n753_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n766_), .A2(KEYINPUT107), .A3(G99gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT107), .B1(new_n766_), .B2(G99gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n765_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n758_), .A2(G106gat), .A3(new_n609_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n752_), .A2(new_n610_), .A3(new_n753_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(G106gat), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n776_), .B(new_n783_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1339gat));
  NAND3_X1  g584(.A1(new_n611_), .A2(new_n612_), .A3(new_n602_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n352_), .A2(new_n787_), .A3(new_n628_), .A4(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n726_), .A2(new_n628_), .A3(new_n664_), .A4(new_n625_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n788_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT111), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n355_), .B(new_n354_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n371_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n346_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n342_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n333_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n801_), .B1(new_n342_), .B2(new_n800_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n329_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n806_), .B2(KEYINPUT56), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n808_), .B(new_n329_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n270_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n347_), .A2(new_n798_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n346_), .A2(KEYINPUT113), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n806_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n373_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT113), .B(new_n329_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(KEYINPUT114), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n623_), .A2(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n814_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n822_), .B2(new_n623_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n324_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n786_), .B1(new_n794_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n325_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n325_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n794_), .A3(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n830_), .A2(new_n837_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT117), .B(G113gat), .Z(new_n839_));
  NAND2_X1  g638(.A1(new_n373_), .A2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT118), .ZN(new_n841_));
  AOI21_X1  g640(.A(G113gat), .B1(new_n828_), .B2(new_n373_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n842_), .A2(KEYINPUT115), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(KEYINPUT115), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n838_), .A2(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(G1340gat));
  NAND3_X1  g644(.A1(new_n830_), .A2(new_n837_), .A3(new_n351_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT119), .B(G120gat), .Z(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n625_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(KEYINPUT60), .B2(new_n847_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n849_), .B1(new_n829_), .B2(new_n851_), .ZN(G1341gat));
  INV_X1    g651(.A(new_n324_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n830_), .A2(new_n837_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G127gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n794_), .A2(new_n827_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n325_), .A2(G127gat), .A3(new_n786_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(G1342gat));
  NAND2_X1  g658(.A1(new_n270_), .A2(G134gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n829_), .B2(new_n623_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(new_n862_), .C1(new_n829_), .C2(new_n623_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n838_), .A2(new_n861_), .B1(new_n864_), .B2(new_n866_), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n612_), .A2(new_n613_), .A3(new_n601_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n856_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n373_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n625_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(G148gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  NOR2_X1   g674(.A1(new_n869_), .A2(new_n325_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT61), .B(G155gat), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  OR3_X1    g677(.A1(new_n869_), .A2(G162gat), .A3(new_n623_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G162gat), .B1(new_n869_), .B2(new_n726_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n608_), .A2(new_n613_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n882_), .A2(new_n431_), .A3(new_n610_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n835_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n373_), .A3(new_n381_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n612_), .A2(new_n373_), .A3(new_n613_), .A4(new_n608_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n609_), .B1(new_n887_), .B2(KEYINPUT122), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(KEYINPUT122), .B2(new_n887_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n835_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n890_), .B2(G169gat), .ZN(new_n891_));
  AOI211_X1 g690(.A(KEYINPUT62), .B(new_n374_), .C1(new_n835_), .C2(new_n889_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n885_), .B1(new_n891_), .B2(new_n892_), .ZN(G1348gat));
  NAND2_X1  g692(.A1(new_n856_), .A2(new_n883_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n894_), .A2(new_n378_), .A3(new_n625_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n835_), .A2(new_n351_), .A3(new_n883_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n378_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT123), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n899_), .A3(new_n378_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n895_), .B1(new_n898_), .B2(new_n900_), .ZN(G1349gat));
  NOR3_X1   g700(.A1(new_n894_), .A2(KEYINPUT124), .A3(new_n325_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(G183gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT124), .B1(new_n894_), .B2(new_n325_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n324_), .A2(new_n402_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n903_), .A2(new_n904_), .B1(new_n884_), .B2(new_n906_), .ZN(G1350gat));
  NAND2_X1  g706(.A1(new_n268_), .A2(new_n403_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT126), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n884_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n835_), .A2(new_n270_), .A3(new_n883_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n911_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(KEYINPUT125), .B1(new_n911_), .B2(G190gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n912_), .B2(new_n913_), .ZN(G1351gat));
  NOR3_X1   g713(.A1(new_n882_), .A2(new_n612_), .A3(new_n609_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n856_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n373_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT127), .B1(new_n917_), .B2(new_n444_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n444_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n916_), .A2(new_n920_), .A3(G197gat), .A4(new_n373_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n918_), .A2(new_n919_), .A3(new_n921_), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n856_), .A2(new_n915_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n625_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n442_), .ZN(G1353gat));
  NAND2_X1  g724(.A1(new_n916_), .A2(new_n853_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  AND2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n926_), .A2(new_n927_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1354gat));
  NAND3_X1  g730(.A1(new_n916_), .A2(new_n434_), .A3(new_n268_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G218gat), .B1(new_n923_), .B2(new_n726_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1355gat));
endmodule


