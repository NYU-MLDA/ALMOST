//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  OAI21_X1  g000(.A(KEYINPUT71), .B1(G169gat), .B2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR3_X1   g002(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT24), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n203_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT25), .B(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT70), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n208_), .B(new_n211_), .C1(new_n212_), .C2(KEYINPUT70), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n213_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT72), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(G176gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n220_), .A2(new_n223_), .A3(KEYINPUT72), .A4(new_n224_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n227_), .A2(new_n205_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n218_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT74), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT31), .ZN(new_n239_));
  INV_X1    g038(.A(G120gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G113gat), .ZN(new_n241_));
  INV_X1    g040(.A(G113gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G120gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT73), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n241_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n246_));
  OAI21_X1  g045(.A(G127gat), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(G120gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n240_), .A2(G113gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT73), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G127gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n241_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n247_), .A2(G134gat), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(G134gat), .B1(new_n247_), .B2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n239_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G134gat), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n245_), .A2(new_n246_), .A3(G127gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n251_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n247_), .A2(new_n253_), .A3(G134gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT31), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n256_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n238_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n256_), .A2(new_n262_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n263_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n256_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n237_), .A3(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G15gat), .B(G43gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n266_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n236_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n264_), .A2(new_n265_), .A3(new_n238_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n237_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n266_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n235_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G197gat), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n288_));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n286_), .B1(new_n284_), .B2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT81), .B1(new_n283_), .B2(G197gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT21), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n287_), .A2(KEYINPUT21), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n289_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n216_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n215_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n221_), .A2(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G183gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT84), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n209_), .A2(G190gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT84), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n302_), .A2(new_n304_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n210_), .A2(new_n313_), .A3(KEYINPUT85), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n306_), .A2(new_n310_), .A3(new_n312_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n207_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT86), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n318_), .A3(new_n207_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n301_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n205_), .B(KEYINPUT87), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n230_), .A2(new_n321_), .A3(new_n225_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n298_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT88), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT20), .B1(new_n298_), .B2(new_n233_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(KEYINPUT83), .B(KEYINPUT20), .C1(new_n298_), .C2(new_n233_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n301_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n315_), .A2(new_n318_), .A3(new_n207_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n318_), .B1(new_n315_), .B2(new_n207_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n322_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n298_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n325_), .A2(new_n328_), .A3(new_n333_), .A4(new_n340_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n290_), .A2(new_n294_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n342_), .A3(new_n322_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n298_), .B2(new_n233_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n327_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G64gat), .B(G92gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT92), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n348_), .A2(KEYINPUT92), .A3(new_n353_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n343_), .A2(new_n328_), .A3(new_n345_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n325_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(new_n327_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n353_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n358_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(new_n357_), .A3(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n362_), .A2(new_n363_), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n353_), .B(new_n360_), .C1(new_n361_), .C2(new_n327_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n358_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n370_));
  INV_X1    g169(.A(G155gat), .ZN(new_n371_));
  INV_X1    g170(.A(G162gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n373_), .A2(KEYINPUT79), .A3(new_n374_), .A4(new_n375_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380_));
  INV_X1    g179(.A(G141gat), .ZN(new_n381_));
  INV_X1    g180(.A(G148gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT3), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT3), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n380_), .A2(new_n385_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT78), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n378_), .B(new_n379_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G141gat), .B(G148gat), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n374_), .A2(KEYINPUT1), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT76), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n373_), .B(new_n375_), .C1(KEYINPUT1), .C2(new_n374_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n392_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n260_), .A2(new_n391_), .A3(new_n396_), .A4(new_n261_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT4), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n397_), .B(new_n401_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n369_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT0), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(G57gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G85gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n369_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n404_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n408_), .B1(new_n403_), .B2(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n397_), .A2(KEYINPUT29), .ZN(new_n416_));
  XOR2_X1   g215(.A(G22gat), .B(G50gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT28), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n416_), .B(new_n418_), .Z(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT80), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(KEYINPUT80), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n397_), .A2(KEYINPUT29), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n298_), .ZN(new_n425_));
  INV_X1    g224(.A(G228gat), .ZN(new_n426_));
  INV_X1    g225(.A(G233gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n342_), .B1(new_n397_), .B2(KEYINPUT29), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n423_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n431_), .A3(new_n423_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AOI211_X1 g234(.A(KEYINPUT82), .B(new_n423_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n420_), .B(new_n421_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n432_), .A2(new_n419_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n434_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n415_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n365_), .A2(new_n368_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n348_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT91), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n362_), .A2(new_n443_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n348_), .A2(KEYINPUT91), .A3(new_n444_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n339_), .B1(new_n338_), .B2(new_n298_), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT88), .B(new_n342_), .C1(new_n337_), .C2(new_n322_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n328_), .B1(new_n453_), .B2(new_n333_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n353_), .B1(new_n454_), .B2(new_n360_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT90), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n414_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n361_), .A2(new_n327_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n363_), .A3(new_n359_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n400_), .A2(new_n369_), .A3(new_n402_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n398_), .A2(new_n410_), .A3(new_n399_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(new_n409_), .A3(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n408_), .B(new_n457_), .C1(new_n403_), .C2(new_n411_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n455_), .A2(new_n460_), .A3(new_n462_), .A4(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n442_), .B1(new_n450_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n282_), .B1(new_n441_), .B2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n413_), .A2(new_n414_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n276_), .A2(new_n281_), .A3(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n437_), .A2(new_n439_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n365_), .A2(new_n472_), .A3(new_n473_), .A4(new_n368_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n474_), .A2(KEYINPUT93), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(KEYINPUT93), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n470_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G230gat), .A2(G233gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT6), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  OR3_X1    g280(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G85gat), .B(G92gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT8), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT10), .B(G99gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n491_), .A2(KEYINPUT64), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(KEYINPUT64), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT66), .B(G92gat), .Z(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(KEYINPUT9), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT65), .B(G85gat), .Z(new_n497_));
  NAND2_X1  g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n496_), .A2(new_n497_), .B1(KEYINPUT9), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n480_), .B(new_n494_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n489_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G71gat), .B(G78gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(KEYINPUT11), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n489_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n478_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(KEYINPUT12), .A3(new_n510_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT12), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n502_), .A2(new_n513_), .A3(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n515_), .B2(new_n478_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n283_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT5), .B(G176gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n516_), .A2(new_n520_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT13), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT13), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT15), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532_));
  INV_X1    g331(.A(G1gat), .ZN(new_n533_));
  INV_X1    g332(.A(G8gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT14), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G8gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n530_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n539_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT69), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n538_), .B(new_n541_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(G229gat), .A3(G233gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(KEYINPUT69), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G169gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n285_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n548_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT16), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n221_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G211gat), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n559_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n538_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n508_), .ZN(new_n564_));
  OR3_X1    g363(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n527_), .A2(new_n554_), .A3(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n477_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n502_), .A2(new_n531_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT67), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT34), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT35), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n574_), .A2(KEYINPUT35), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n571_), .B(new_n579_), .C1(new_n502_), .C2(new_n541_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n576_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT36), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n585_), .A2(KEYINPUT36), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n582_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n570_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n587_), .B(KEYINPUT37), .C1(new_n582_), .C2(new_n590_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n569_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n569_), .A2(KEYINPUT94), .A3(new_n594_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n471_), .A2(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT95), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(KEYINPUT95), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(KEYINPUT38), .A3(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n588_), .A2(new_n591_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n569_), .A2(new_n415_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(G1gat), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT38), .B1(new_n601_), .B2(new_n602_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1324gat));
  NAND2_X1  g409(.A1(new_n365_), .A2(new_n368_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n569_), .A2(new_n611_), .A3(new_n605_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G8gat), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT96), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n597_), .A2(new_n534_), .A3(new_n611_), .A4(new_n598_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n613_), .A2(KEYINPUT96), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n614_), .A2(new_n619_), .A3(new_n615_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT98), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n618_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(new_n282_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n569_), .A2(new_n627_), .A3(new_n605_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(G15gat), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n629_), .B1(new_n628_), .B2(G15gat), .ZN(new_n633_));
  OR3_X1    g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n282_), .A2(G15gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n597_), .A2(new_n598_), .A3(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n635_), .A3(new_n637_), .ZN(G1326gat));
  XNOR2_X1  g437(.A(new_n442_), .B(KEYINPUT100), .ZN(new_n639_));
  INV_X1    g438(.A(G22gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT101), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n597_), .A2(new_n598_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n569_), .A2(new_n605_), .A3(new_n639_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(G22gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n644_), .B2(G22gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT102), .Z(G1327gat));
  NAND4_X1  g448(.A1(new_n525_), .A2(new_n526_), .A3(new_n553_), .A4(new_n567_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT103), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n462_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n455_), .A2(new_n462_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n652_), .A2(new_n356_), .B1(new_n653_), .B2(new_n358_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT93), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n473_), .A4(new_n472_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n474_), .A2(KEYINPUT93), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT43), .B(new_n594_), .C1(new_n658_), .C2(new_n470_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n592_), .A2(new_n593_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n477_), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n651_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT44), .B(new_n651_), .C1(new_n659_), .C2(new_n662_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n665_), .A2(G29gat), .A3(new_n415_), .A4(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n477_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n605_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n650_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(new_n471_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(G29gat), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT104), .ZN(G1328gat));
  NAND3_X1  g473(.A1(new_n665_), .A2(new_n611_), .A3(new_n666_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n665_), .A2(new_n677_), .A3(new_n611_), .A4(new_n666_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(G36gat), .A3(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n671_), .A2(G36gat), .A3(new_n654_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(KEYINPUT46), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n665_), .A2(new_n627_), .A3(new_n666_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G43gat), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n671_), .A2(G43gat), .A3(new_n282_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g491(.A(new_n671_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G50gat), .B1(new_n693_), .B2(new_n639_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n665_), .A2(new_n666_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n442_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(G1331gat));
  INV_X1    g496(.A(new_n567_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n527_), .A2(new_n554_), .A3(new_n698_), .A4(new_n605_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n668_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(G57gat), .A3(new_n415_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(new_n702_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n525_), .A2(new_n526_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n594_), .A2(new_n554_), .A3(new_n698_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n668_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n415_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n703_), .A2(new_n704_), .A3(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n611_), .A2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT109), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n700_), .A2(new_n611_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G64gat), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT108), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(new_n717_), .A3(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT48), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n714_), .B2(G64gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT108), .B(new_n710_), .C1(new_n700_), .C2(new_n611_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n713_), .B1(new_n719_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT110), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n707_), .A2(new_n726_), .A3(new_n627_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n700_), .A2(new_n627_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G71gat), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT49), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT49), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n707_), .A2(new_n733_), .A3(new_n639_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n700_), .A2(new_n639_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G78gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n737_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n738_), .B2(new_n739_), .ZN(G1335gat));
  NAND3_X1  g539(.A1(new_n527_), .A2(new_n554_), .A3(new_n567_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n668_), .A2(new_n605_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n415_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n659_), .A2(new_n662_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n741_), .B(KEYINPUT112), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n415_), .A2(new_n497_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n742_), .B2(new_n611_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n654_), .A2(new_n495_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT113), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n747_), .B2(new_n752_), .ZN(G1337gat));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  INV_X1    g553(.A(G99gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n747_), .B2(new_n627_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n492_), .A2(new_n493_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n742_), .A2(new_n627_), .A3(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n754_), .B1(new_n760_), .B2(KEYINPUT51), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n759_), .A2(KEYINPUT114), .A3(new_n762_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n759_), .A2(KEYINPUT115), .A3(new_n762_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT115), .B1(new_n759_), .B2(new_n762_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n761_), .A2(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n742_), .A2(new_n490_), .A3(new_n442_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n747_), .A2(new_n442_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(G106gat), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT52), .B(new_n490_), .C1(new_n747_), .C2(new_n442_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n767_), .B(new_n774_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n611_), .A2(new_n442_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n282_), .A2(new_n471_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780_));
  INV_X1    g579(.A(new_n478_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n512_), .A2(new_n781_), .A3(new_n514_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n510_), .A2(KEYINPUT12), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n507_), .B1(new_n489_), .B2(new_n501_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n514_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n478_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n515_), .A2(new_n790_), .A3(new_n478_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n783_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n520_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n548_), .A2(new_n552_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n539_), .A2(G229gat), .A3(G233gat), .A4(new_n542_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n551_), .B1(new_n545_), .B2(new_n540_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n790_), .B1(new_n515_), .B2(new_n478_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT55), .B(new_n781_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n782_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n520_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n793_), .A2(new_n521_), .A3(new_n797_), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n661_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n780_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n804_), .A2(new_n805_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT117), .A3(new_n661_), .A4(new_n806_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n793_), .A2(new_n521_), .A3(new_n553_), .A4(new_n803_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n797_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n604_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT116), .B1(new_n814_), .B2(KEYINPUT57), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(new_n811_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(KEYINPUT116), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n812_), .A2(new_n813_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n605_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(KEYINPUT57), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n567_), .B1(new_n816_), .B2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n706_), .A2(new_n527_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n706_), .A2(KEYINPUT54), .A3(new_n527_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n779_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n553_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n824_), .A2(new_n829_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n779_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n833_), .B2(KEYINPUT118), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(KEYINPUT118), .B2(new_n833_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n821_), .A2(new_n822_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n810_), .A2(new_n661_), .A3(new_n806_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n698_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n827_), .A2(new_n828_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n835_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n553_), .A2(G113gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT119), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n831_), .B1(new_n845_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n844_), .B2(new_n705_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n835_), .A2(KEYINPUT121), .A3(new_n527_), .A4(new_n843_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(G120gat), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT60), .ZN(new_n853_));
  AOI21_X1  g652(.A(G120gat), .B1(new_n527_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n853_), .B2(G120gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n830_), .A2(new_n856_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n852_), .A2(new_n859_), .ZN(G1341gat));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n567_), .B2(new_n251_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n843_), .B(new_n862_), .C1(new_n830_), .C2(new_n836_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G127gat), .B1(new_n863_), .B2(KEYINPUT122), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n698_), .A3(new_n830_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(KEYINPUT123), .A3(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1342gat));
  OAI21_X1  g669(.A(G134gat), .B1(new_n844_), .B2(new_n594_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n830_), .A2(new_n257_), .A3(new_n604_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1343gat));
  AOI21_X1  g672(.A(new_n627_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n611_), .A2(new_n473_), .A3(new_n471_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n554_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n381_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n705_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n382_), .ZN(G1345gat));
  OR3_X1    g679(.A1(new_n876_), .A2(KEYINPUT124), .A3(new_n567_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT124), .B1(new_n876_), .B2(new_n567_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT61), .B(G155gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(new_n884_), .A3(new_n882_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n876_), .B2(new_n594_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n604_), .A2(new_n372_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n876_), .B2(new_n890_), .ZN(G1347gat));
  OR2_X1    g690(.A1(new_n841_), .A2(new_n842_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n611_), .A2(new_n472_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n639_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895_), .B2(new_n554_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n228_), .A3(new_n553_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n897_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n900_), .A3(new_n901_), .ZN(G1348gat));
  AOI21_X1  g701(.A(G176gat), .B1(new_n899_), .B2(new_n527_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n442_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n705_), .A2(new_n229_), .A3(new_n893_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1349gat));
  NOR2_X1   g705(.A1(new_n893_), .A2(new_n567_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(KEYINPUT125), .A3(new_n907_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n221_), .A3(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n567_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n899_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n917_), .A3(new_n914_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n895_), .B2(new_n594_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n604_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n895_), .B2(new_n921_), .ZN(G1351gat));
  AND2_X1   g721(.A1(new_n611_), .A2(new_n440_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n874_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n554_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n285_), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n705_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n283_), .ZN(G1353gat));
  AOI21_X1  g727(.A(new_n567_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n874_), .A2(new_n923_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT127), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n874_), .A2(new_n932_), .A3(new_n923_), .A4(new_n929_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n924_), .B2(new_n594_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n605_), .A2(G218gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n924_), .B2(new_n938_), .ZN(G1355gat));
endmodule


