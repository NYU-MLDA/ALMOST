//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  INV_X1    g004(.A(G141gat), .ZN(new_n206_));
  INV_X1    g005(.A(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n219_));
  AND2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n220_), .A2(KEYINPUT1), .B1(new_n206_), .B2(new_n207_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n222_), .A3(new_n216_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n223_), .A3(new_n209_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n218_), .A2(new_n219_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n219_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n204_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT95), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n224_), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n204_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT95), .B(new_n204_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n229_), .A2(KEYINPUT4), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n234_), .B(new_n204_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT96), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(KEYINPUT89), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n218_), .A2(new_n224_), .A3(new_n219_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n240_), .A2(KEYINPUT96), .A3(new_n234_), .A4(new_n204_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n244_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G85gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G57gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n252_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n248_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n244_), .B1(new_n233_), .B2(new_n242_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT101), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT101), .B(new_n254_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n263_), .A2(G204gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT90), .B(G204gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(G197gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n262_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G197gat), .A2(G204gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n265_), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT21), .B(new_n269_), .C1(new_n270_), .C2(G197gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n262_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n266_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  INV_X1    g076(.A(G169gat), .ZN(new_n278_));
  INV_X1    g077(.A(G176gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT25), .B(G183gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n288_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n288_), .B2(new_n292_), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT23), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G183gat), .A3(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n293_), .A2(new_n294_), .A3(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(KEYINPUT22), .B(G169gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT85), .B(G176gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n283_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n300_), .B1(G183gat), .B2(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n276_), .B1(new_n304_), .B2(new_n312_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n268_), .A2(new_n271_), .B1(new_n274_), .B2(KEYINPUT21), .ZN(new_n314_));
  AND2_X1   g113(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n296_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n300_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n309_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n280_), .A2(new_n301_), .A3(new_n281_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n321_), .A2(new_n300_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n281_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT84), .B(new_n323_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT84), .B1(new_n282_), .B2(new_n323_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n322_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n295_), .B2(KEYINPUT25), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT81), .A3(G183gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT25), .B1(new_n315_), .B2(new_n316_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n290_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT82), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n334_), .A2(new_n335_), .A3(new_n338_), .A4(new_n290_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n314_), .B(new_n320_), .C1(new_n329_), .C2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n313_), .A2(KEYINPUT20), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G226gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT19), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n320_), .B1(new_n340_), .B2(new_n329_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n276_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n288_), .A2(new_n292_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT92), .ZN(new_n349_));
  INV_X1    g148(.A(new_n303_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n288_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n314_), .A3(new_n311_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n344_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n347_), .A2(new_n353_), .A3(KEYINPUT20), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT93), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n346_), .B2(new_n276_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT93), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n354_), .A4(new_n353_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n345_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G92gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT18), .B(G64gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n345_), .A2(new_n356_), .A3(new_n365_), .A4(new_n360_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n230_), .A2(KEYINPUT29), .ZN(new_n373_));
  OAI211_X1 g172(.A(G228gat), .B(G233gat), .C1(new_n314_), .C2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT29), .B1(new_n225_), .B2(new_n226_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n276_), .ZN(new_n377_));
  INV_X1    g176(.A(G22gat), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n372_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OR4_X1    g180(.A1(KEYINPUT28), .A2(new_n225_), .A3(new_n226_), .A4(KEYINPUT29), .ZN(new_n382_));
  INV_X1    g181(.A(G50gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT28), .B1(new_n240_), .B2(KEYINPUT29), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n374_), .A2(new_n377_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G22gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n372_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n381_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n387_), .B1(new_n381_), .B2(new_n392_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n342_), .A2(new_n344_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n354_), .B1(new_n358_), .B2(new_n353_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n368_), .B(KEYINPUT27), .C1(new_n398_), .C2(new_n365_), .ZN(new_n399_));
  AND4_X1   g198(.A1(new_n261_), .A2(new_n371_), .A3(new_n395_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n398_), .B(new_n402_), .C1(new_n361_), .C2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n401_), .B1(new_n361_), .B2(KEYINPUT100), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n260_), .A3(new_n259_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT94), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n369_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n367_), .A2(KEYINPUT94), .A3(new_n368_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n252_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT97), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT33), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n257_), .A2(KEYINPUT97), .A3(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n233_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n417_), .A2(KEYINPUT99), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(KEYINPUT99), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n252_), .B1(new_n247_), .B2(new_n244_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT98), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT98), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n422_), .B(new_n252_), .C1(new_n247_), .C2(new_n244_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n416_), .A3(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n407_), .B1(new_n411_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n395_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n400_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(G43gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(G43gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n430_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n442_), .A2(KEYINPUT88), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n438_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT86), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n430_), .A2(KEYINPUT87), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n430_), .A2(KEYINPUT87), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n442_), .A2(KEYINPUT88), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n443_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT102), .B1(new_n428_), .B2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n371_), .A2(new_n399_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n453_), .A2(new_n261_), .A3(new_n427_), .A4(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT102), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n443_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n257_), .A2(KEYINPUT97), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n421_), .A2(new_n423_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n417_), .B(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(KEYINPUT33), .A2(new_n459_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n463_), .A2(new_n416_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n395_), .B1(new_n464_), .B2(new_n407_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n457_), .B(new_n458_), .C1(new_n465_), .C2(new_n400_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n454_), .A2(new_n456_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G85gat), .B(G92gat), .Z(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(KEYINPUT9), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT10), .B(G99gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT64), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n478_), .B2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(KEYINPUT9), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT7), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n472_), .B(new_n473_), .C1(new_n483_), .C2(KEYINPUT7), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n475_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT8), .B1(new_n475_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  OAI221_X1 g290(.A(new_n475_), .B1(new_n489_), .B2(KEYINPUT8), .C1(new_n486_), .C2(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n482_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G29gat), .B(G36gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G43gat), .B(G50gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n469_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  OAI221_X1 g297(.A(new_n476_), .B1(KEYINPUT9), .B2(new_n480_), .C1(new_n478_), .C2(G106gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(KEYINPUT15), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G232gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n498_), .B(new_n502_), .C1(KEYINPUT35), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(KEYINPUT35), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(KEYINPUT36), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n468_), .B1(new_n509_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(KEYINPUT71), .A3(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(KEYINPUT36), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(new_n515_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(KEYINPUT37), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT72), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n522_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n523_), .A2(new_n524_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n525_), .B2(KEYINPUT37), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n467_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n531_));
  XOR2_X1   g330(.A(G71gat), .B(G78gat), .Z(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n482_), .B2(new_n493_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n499_), .A2(new_n535_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n500_), .B2(KEYINPUT67), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  INV_X1    g342(.A(new_n493_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n499_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n537_), .B1(new_n545_), .B2(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT68), .B(G204gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT5), .B(G176gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n555_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G15gat), .B(G22gat), .Z(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT73), .B(G1gat), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G8gat), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n566_), .B2(KEYINPUT14), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G1gat), .B(G8gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n497_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT76), .ZN(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n497_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n571_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT77), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(new_n570_), .A3(KEYINPUT76), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n572_), .A2(new_n501_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n577_), .A3(new_n570_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT79), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n263_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT78), .B(G169gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(KEYINPUT79), .A3(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n563_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n569_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n536_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n543_), .A3(KEYINPUT17), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n600_), .A2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n600_), .B(new_n606_), .C1(KEYINPUT17), .C2(new_n605_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT75), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n528_), .A2(new_n597_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n565_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n261_), .B(KEYINPUT103), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT38), .ZN(new_n616_));
  INV_X1    g415(.A(new_n609_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n597_), .B(KEYINPUT104), .ZN(new_n618_));
  INV_X1    g417(.A(new_n525_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n467_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT105), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(KEYINPUT105), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n617_), .B(new_n618_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n261_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n616_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT106), .Z(G1324gat));
  INV_X1    g425(.A(G8gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n455_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n612_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G8gat), .B1(new_n623_), .B2(new_n455_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT107), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT107), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n633_), .B(G8gat), .C1(new_n623_), .C2(new_n455_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n631_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n632_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n629_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT40), .B(new_n629_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n623_), .B2(new_n458_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  INV_X1    g442(.A(G15gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n612_), .A2(new_n644_), .A3(new_n453_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1326gat));
  OAI21_X1  g445(.A(G22gat), .B1(new_n623_), .B2(new_n427_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT42), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n395_), .A2(new_n378_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT108), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n612_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(G1327gat));
  AND3_X1   g451(.A1(new_n467_), .A2(new_n525_), .A3(new_n610_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n597_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT112), .ZN(new_n655_));
  INV_X1    g454(.A(new_n261_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n614_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT111), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n467_), .A2(new_n526_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(KEYINPUT43), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT109), .B(new_n663_), .C1(new_n467_), .C2(new_n526_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n467_), .A2(new_n663_), .A3(new_n526_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n662_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n618_), .A2(new_n610_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n659_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n661_), .A2(KEYINPUT43), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT109), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n661_), .A2(new_n660_), .A3(KEYINPUT43), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n665_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n668_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n670_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n669_), .B(KEYINPUT44), .C1(new_n676_), .C2(new_n659_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n662_), .A2(new_n664_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n668_), .B1(new_n679_), .B2(new_n665_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT111), .B(new_n678_), .C1(new_n680_), .C2(new_n670_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n658_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n657_), .B1(new_n682_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n669_), .A2(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n674_), .A2(new_n675_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n659_), .B1(new_n687_), .B2(KEYINPUT110), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n681_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n685_), .B1(new_n689_), .B2(new_n628_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n655_), .A2(new_n685_), .A3(new_n628_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n684_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n455_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n695_), .B(KEYINPUT46), .C1(new_n696_), .C2(new_n685_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n697_), .ZN(G1329gat));
  INV_X1    g497(.A(G43gat), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n699_), .B(new_n458_), .C1(new_n677_), .C2(new_n681_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n655_), .A2(new_n453_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT47), .B1(new_n700_), .B2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n689_), .A2(G43gat), .A3(new_n453_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n704_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1330gat));
  NAND3_X1  g509(.A1(new_n655_), .A2(new_n383_), .A3(new_n395_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n689_), .A2(new_n395_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT114), .B1(new_n712_), .B2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n427_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT114), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n383_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n713_), .B2(new_n716_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n563_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n596_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n610_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n528_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n614_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n621_), .A2(new_n622_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n720_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n656_), .A2(G57gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n725_), .B2(new_n455_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT48), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n455_), .A2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n721_), .B2(new_n731_), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n725_), .B2(new_n458_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT49), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n458_), .A2(G71gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT115), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n721_), .B2(new_n736_), .ZN(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n725_), .B2(new_n427_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT50), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n721_), .A2(G78gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n427_), .B2(new_n740_), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n718_), .A2(new_n719_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n674_), .A2(new_n610_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(G85gat), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n261_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n653_), .A2(new_n614_), .A3(new_n742_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(new_n746_), .ZN(G1336gat));
  INV_X1    g546(.A(G92gat), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n743_), .A2(new_n748_), .A3(new_n455_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n653_), .A2(new_n628_), .A3(new_n742_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(new_n750_), .ZN(G1337gat));
  NAND2_X1  g550(.A1(new_n653_), .A2(new_n742_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n752_), .A2(new_n458_), .A3(new_n478_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G99gat), .B1(new_n743_), .B2(new_n458_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT117), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n756_), .A3(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n758_), .A2(KEYINPUT118), .A3(KEYINPUT51), .A4(new_n760_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n758_), .A2(KEYINPUT51), .A3(new_n760_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT118), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n762_), .B2(new_n765_), .ZN(G1338gat));
  OR3_X1    g565(.A1(new_n752_), .A2(G106gat), .A3(new_n427_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G106gat), .B1(new_n743_), .B2(new_n427_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT52), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT53), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n767_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1339gat));
  NOR2_X1   g574(.A1(new_n458_), .A2(new_n395_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(new_n628_), .A3(new_n658_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n575_), .A2(new_n578_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n577_), .B1(new_n583_), .B2(new_n570_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n593_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n579_), .A2(new_n586_), .A3(new_n592_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n559_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT121), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n548_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n539_), .A2(new_n541_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n537_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n541_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n549_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n792_), .B2(KEYINPUT55), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n547_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(KEYINPUT120), .A3(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n787_), .B1(new_n793_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n555_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n792_), .A2(new_n788_), .A3(KEYINPUT55), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT120), .B1(new_n794_), .B2(new_n795_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n548_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n798_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n797_), .A2(new_n801_), .A3(KEYINPUT56), .A4(new_n798_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n719_), .A3(new_n556_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n525_), .B1(new_n786_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT124), .A3(KEYINPUT57), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n596_), .B(new_n557_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT57), .B(new_n619_), .C1(new_n810_), .C2(new_n785_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n782_), .A2(new_n783_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n805_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n804_), .A2(KEYINPUT122), .A3(new_n805_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n556_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT58), .A4(new_n556_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n526_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT123), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n808_), .A2(KEYINPUT57), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n822_), .A2(new_n526_), .A3(new_n827_), .A4(new_n823_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n814_), .A2(new_n825_), .A3(new_n826_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT125), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n813_), .A2(new_n809_), .B1(new_n824_), .B2(KEYINPUT123), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n826_), .A4(new_n828_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(new_n833_), .A3(new_n609_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n527_), .A2(new_n596_), .A3(new_n718_), .A4(new_n611_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n779_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n719_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n837_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n778_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n814_), .A2(new_n826_), .A3(new_n824_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n610_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(new_n837_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n845_), .A2(KEYINPUT59), .A3(new_n779_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n719_), .A2(G113gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n839_), .B1(new_n847_), .B2(new_n848_), .ZN(G1340gat));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n846_), .B(new_n563_), .C1(new_n850_), .C2(new_n838_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n718_), .B2(G120gat), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n838_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G120gat), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g656(.A(G127gat), .B1(new_n838_), .B2(new_n611_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n617_), .A2(G127gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n847_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n841_), .B2(new_n619_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(KEYINPUT126), .B(new_n861_), .C1(new_n841_), .C2(new_n619_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n527_), .A2(new_n861_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n842_), .A2(new_n846_), .A3(new_n866_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n864_), .A2(new_n865_), .A3(new_n867_), .ZN(G1343gat));
  AOI21_X1  g667(.A(new_n658_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n453_), .A2(new_n427_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n628_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n596_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n206_), .ZN(G1344gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n718_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n207_), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n873_), .A2(new_n610_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n873_), .A2(new_n881_), .A3(new_n527_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n873_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n525_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n881_), .B2(new_n884_), .ZN(G1347gat));
  NOR3_X1   g684(.A1(new_n777_), .A2(new_n455_), .A3(new_n614_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n845_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n278_), .B1(new_n888_), .B2(new_n719_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n845_), .A2(new_n305_), .A3(new_n596_), .A4(new_n887_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT62), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(KEYINPUT62), .B2(new_n889_), .ZN(G1348gat));
  AOI21_X1  g691(.A(new_n306_), .B1(new_n888_), .B2(new_n563_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n887_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n718_), .A2(new_n279_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n611_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n609_), .A2(new_n291_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n897_), .A2(new_n317_), .B1(new_n888_), .B2(new_n898_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n888_), .A2(new_n290_), .A3(new_n525_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n845_), .A2(new_n527_), .A3(new_n887_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n296_), .B2(new_n901_), .ZN(G1351gat));
  AOI21_X1  g701(.A(new_n871_), .B1(new_n834_), .B2(new_n837_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n455_), .A2(new_n656_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n719_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G197gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n263_), .A3(new_n719_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1352gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n563_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G204gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n270_), .B2(new_n910_), .ZN(G1353gat));
  NAND3_X1  g711(.A1(new_n903_), .A2(new_n617_), .A3(new_n904_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  NAND4_X1  g716(.A1(new_n840_), .A2(new_n525_), .A3(new_n870_), .A4(new_n904_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT127), .ZN(new_n919_));
  INV_X1    g718(.A(G218gat), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n903_), .A2(new_n921_), .A3(new_n525_), .A4(new_n904_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n920_), .A3(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n905_), .A2(G218gat), .A3(new_n526_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1355gat));
endmodule


