//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n208_), .B(new_n211_), .Z(new_n212_));
  NAND2_X1  g011(.A1(G229gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(new_n208_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n208_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n214_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n212_), .A2(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G113gat), .B(G141gat), .Z(new_n220_));
  XNOR2_X1  g019(.A(G169gat), .B(G197gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n219_), .A2(new_n222_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT79), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G85gat), .ZN(new_n233_));
  INV_X1    g032(.A(G92gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n229_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  NOR4_X1   g037(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT6), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(G99gat), .B2(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n248_));
  OAI22_X1  g047(.A1(new_n246_), .A2(new_n248_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n238_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT8), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n235_), .A2(KEYINPUT9), .A3(new_n229_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI22_X1  g057(.A1(new_n246_), .A2(new_n248_), .B1(KEYINPUT9), .B2(new_n229_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT64), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n245_), .A2(G99gat), .A3(G106gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT9), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n261_), .A2(new_n262_), .B1(new_n230_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n256_), .A4(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n238_), .B(KEYINPUT8), .C1(new_n244_), .C2(new_n249_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n252_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT67), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n252_), .A2(new_n267_), .A3(new_n271_), .A4(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n275_));
  XOR2_X1   g074(.A(G71gat), .B(G78gat), .Z(new_n276_));
  AND2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(KEYINPUT11), .B2(new_n274_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n275_), .A2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT12), .B1(new_n273_), .B2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n270_), .A2(new_n272_), .A3(new_n280_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n269_), .A3(KEYINPUT12), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G230gat), .ZN(new_n287_));
  INV_X1    g086(.A(G233gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n273_), .A2(new_n281_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n292_), .B2(new_n283_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n294_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G120gat), .B(G148gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(G176gat), .B(G204gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT70), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n303_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT13), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n296_), .A2(new_n297_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(new_n304_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n314_), .B2(new_n307_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n228_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G155gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT16), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n208_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(new_n280_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n321_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT17), .B1(new_n324_), .B2(new_n321_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT17), .B(new_n321_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n316_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT103), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n316_), .A2(KEYINPUT103), .A3(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G232gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT34), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n270_), .A2(new_n211_), .A3(new_n272_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n270_), .A2(KEYINPUT73), .A3(new_n211_), .A4(new_n272_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n269_), .A2(new_n215_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n341_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  AOI211_X1 g148(.A(new_n340_), .B(new_n349_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G134gat), .B(G162gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G190gat), .B(G218gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT75), .Z(new_n356_));
  NOR3_X1   g155(.A1(new_n348_), .A2(new_n350_), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n353_), .B(KEYINPUT36), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(KEYINPUT76), .B(new_n358_), .C1(new_n348_), .C2(new_n350_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n357_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G183gat), .A3(G190gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n368_), .A3(KEYINPUT84), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n365_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371_));
  INV_X1    g170(.A(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n369_), .B(new_n370_), .C1(G183gat), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G169gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT22), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT22), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G169gat), .ZN(new_n380_));
  INV_X1    g179(.A(G176gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n382_), .B2(KEYINPUT83), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n376_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT81), .B1(new_n372_), .B2(KEYINPUT26), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n373_), .A2(KEYINPUT26), .A3(new_n374_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT25), .B(G183gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n366_), .A2(new_n368_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT24), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n400_), .B1(new_n385_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n392_), .A2(new_n393_), .A3(KEYINPUT82), .A4(new_n394_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n387_), .B1(new_n397_), .B2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G71gat), .B(G99gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G43gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n406_), .B(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT31), .Z(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT86), .B(G15gat), .Z(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(KEYINPUT85), .B(KEYINPUT30), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G113gat), .B(G120gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G134gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G127gat), .ZN(new_n419_));
  INV_X1    g218(.A(G127gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G134gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n417_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n420_), .A2(G134gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n418_), .A2(G127gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT87), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n416_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n415_), .B(new_n431_), .Z(new_n432_));
  OR2_X1    g231(.A1(new_n410_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n410_), .A2(new_n432_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G155gat), .A2(G162gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n436_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT89), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(KEYINPUT90), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G141gat), .A2(G148gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT2), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT2), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(G141gat), .A3(G148gat), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n442_), .A2(new_n445_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT89), .B1(new_n443_), .B2(KEYINPUT90), .ZN(new_n451_));
  NOR3_X1   g250(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(KEYINPUT90), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n440_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n442_), .A2(new_n446_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT1), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n436_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458_));
  INV_X1    g257(.A(G155gat), .ZN(new_n459_));
  INV_X1    g258(.A(G162gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n437_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n455_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n454_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT28), .Z(new_n467_));
  INV_X1    g266(.A(G218gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G211gat), .ZN(new_n469_));
  INV_X1    g268(.A(G211gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G218gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n473_));
  INV_X1    g272(.A(G197gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G204gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT21), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(G197gat), .B2(G204gat), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n472_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(G204gat), .A3(new_n477_), .ZN(new_n482_));
  OR3_X1    g281(.A1(new_n474_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT92), .B1(new_n474_), .B2(G204gat), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n479_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n479_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n467_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n466_), .B(KEYINPUT28), .ZN(new_n493_));
  INV_X1    g292(.A(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G78gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G106gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G22gat), .B(G50gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n492_), .A2(new_n495_), .A3(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n431_), .B1(new_n454_), .B2(new_n463_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n461_), .A2(new_n437_), .B1(G155gat), .B2(G162gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n445_), .A2(new_n442_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n447_), .A2(new_n449_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n444_), .B1(new_n511_), .B2(KEYINPUT3), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n441_), .A2(new_n443_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n457_), .A2(new_n462_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n455_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n515_), .A2(new_n518_), .A3(new_n430_), .A4(new_n425_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(new_n519_), .A3(KEYINPUT4), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n506_), .A2(new_n519_), .A3(KEYINPUT97), .A4(KEYINPUT4), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G225gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n506_), .B2(KEYINPUT4), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n506_), .A2(new_n519_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n530_), .A2(new_n526_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G1gat), .B(G29gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G85gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT0), .B(G57gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT102), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n527_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n536_), .B1(new_n540_), .B2(new_n531_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n539_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n505_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(G183gat), .A2(G190gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n398_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n382_), .A2(new_n384_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n382_), .A2(KEYINPUT94), .A3(new_n384_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n402_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G190gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n394_), .A2(new_n553_), .ZN(new_n554_));
  AND4_X1   g353(.A1(new_n552_), .A2(new_n554_), .A3(new_n370_), .A4(new_n369_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n490_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n395_), .A2(new_n396_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(new_n404_), .A3(new_n403_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n485_), .A2(new_n481_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(new_n387_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n560_), .A3(KEYINPUT20), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n562_));
  AND2_X1   g361(.A1(G226gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n366_), .A2(new_n368_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(G183gat), .B2(G190gat), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n382_), .A2(KEYINPUT94), .A3(new_n384_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT94), .B1(new_n382_), .B2(new_n384_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n552_), .A2(new_n554_), .A3(new_n370_), .A4(new_n369_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n559_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n564_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n573_), .A2(KEYINPUT20), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n559_), .B1(new_n558_), .B2(new_n387_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT95), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n406_), .A2(new_n490_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT95), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n572_), .A4(new_n574_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n565_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G8gat), .B(G36gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT18), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G64gat), .B(G92gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n565_), .A2(new_n577_), .A3(new_n580_), .A4(new_n585_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT27), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(KEYINPUT96), .A3(new_n586_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n561_), .A2(new_n564_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT100), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT99), .B(KEYINPUT20), .Z(new_n596_));
  AND3_X1   g395(.A1(new_n572_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n572_), .B2(new_n596_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n576_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n594_), .B1(new_n599_), .B2(new_n573_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n586_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(KEYINPUT27), .A3(new_n589_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n593_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n544_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n585_), .A2(KEYINPUT32), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n605_), .B1(new_n581_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n575_), .A2(new_n576_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n609_), .A2(new_n579_), .B1(new_n564_), .B2(new_n561_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n610_), .A2(KEYINPUT98), .A3(new_n577_), .A4(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n538_), .A2(new_n541_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n600_), .A2(new_n607_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n590_), .A2(new_n592_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n536_), .B1(new_n530_), .B2(new_n525_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n506_), .A2(KEYINPUT4), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n526_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n524_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n531_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n623_), .B2(new_n537_), .ZN(new_n624_));
  NOR4_X1   g423(.A1(new_n540_), .A2(KEYINPUT33), .A3(new_n531_), .A4(new_n536_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n615_), .B1(new_n616_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n505_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n604_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n627_), .A2(KEYINPUT101), .A3(new_n628_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n435_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n603_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n628_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n542_), .A2(new_n543_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n435_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n364_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n335_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n636_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G1gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT37), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n357_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n359_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(new_n330_), .C1(new_n363_), .C2(KEYINPUT37), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT78), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT78), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n311_), .A2(new_n315_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n649_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n538_), .A2(KEYINPUT33), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n623_), .A2(new_n622_), .A3(new_n537_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n620_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n590_), .A2(new_n592_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n538_), .A2(new_n541_), .B1(new_n600_), .B2(new_n607_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n656_), .A2(new_n657_), .B1(new_n612_), .B2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n630_), .B1(new_n659_), .B2(new_n505_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n604_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n632_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n435_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n638_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n228_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n653_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n203_), .A3(new_n641_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(KEYINPUT104), .A3(new_n644_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT104), .B1(new_n667_), .B2(new_n644_), .ZN(new_n669_));
  OAI221_X1 g468(.A(new_n643_), .B1(new_n644_), .B2(new_n667_), .C1(new_n668_), .C2(new_n669_), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n335_), .A2(new_n639_), .A3(new_n634_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n204_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n639_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n603_), .A3(new_n333_), .A4(new_n334_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(KEYINPUT106), .A3(G8gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n676_), .A3(KEYINPUT39), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n671_), .B(new_n678_), .C1(new_n672_), .C2(new_n204_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n634_), .A2(G8gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n666_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT105), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n666_), .A2(new_n683_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n677_), .A2(new_n679_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n677_), .A2(new_n685_), .A3(KEYINPUT40), .A4(new_n679_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  INV_X1    g489(.A(G15gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n666_), .A2(new_n691_), .A3(new_n435_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n640_), .A2(new_n435_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n693_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT41), .B1(new_n693_), .B2(G15gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n692_), .B1(new_n694_), .B2(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(G22gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n666_), .A2(new_n697_), .A3(new_n505_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n640_), .A2(new_n505_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n699_), .A2(G22gat), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT108), .B(new_n698_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1327gat));
  INV_X1    g506(.A(new_n330_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n363_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n652_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n665_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G29gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n641_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n316_), .A2(new_n708_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n647_), .B1(new_n363_), .B2(KEYINPUT37), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT109), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n647_), .C1(new_n363_), .C2(KEYINPUT37), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n719_), .B2(new_n664_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n721_), .B(new_n715_), .C1(new_n633_), .C2(new_n638_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n714_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT110), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n715_), .A2(new_n721_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n662_), .A2(new_n663_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n638_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n716_), .B(new_n718_), .C1(new_n633_), .C2(new_n638_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(KEYINPUT43), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n725_), .B(new_n726_), .C1(new_n732_), .C2(new_n714_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n724_), .A2(new_n733_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n726_), .B(new_n714_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n636_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT111), .B1(new_n737_), .B2(G29gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n739_), .B(new_n712_), .C1(new_n734_), .C2(new_n736_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n713_), .B1(new_n738_), .B2(new_n740_), .ZN(G1328gat));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n735_), .A2(new_n634_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n734_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n634_), .A2(G36gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n665_), .A2(new_n710_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT112), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n665_), .A2(new_n749_), .A3(new_n710_), .A4(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n742_), .B1(new_n745_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n751_), .B(KEYINPUT45), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n720_), .A2(new_n722_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n714_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(KEYINPUT44), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n603_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n724_), .B2(new_n733_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n755_), .B(KEYINPUT46), .C1(new_n760_), .C2(new_n743_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n754_), .A2(new_n761_), .ZN(G1329gat));
  NAND2_X1  g561(.A1(new_n435_), .A2(G43gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n735_), .B(new_n763_), .C1(new_n724_), .C2(new_n733_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n711_), .A2(new_n435_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT113), .B(G43gat), .Z(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT47), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n769_));
  INV_X1    g568(.A(new_n767_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n734_), .A2(new_n758_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n769_), .B(new_n770_), .C1(new_n771_), .C2(new_n763_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n768_), .A2(new_n772_), .ZN(G1330gat));
  AOI21_X1  g572(.A(G50gat), .B1(new_n711_), .B2(new_n505_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n771_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n505_), .A2(G50gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(G1331gat));
  INV_X1    g576(.A(G57gat), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n649_), .A2(new_n650_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n228_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n664_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n779_), .A2(new_n781_), .A3(new_n652_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n782_), .B2(new_n636_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT114), .Z(new_n784_));
  NOR2_X1   g583(.A1(new_n780_), .A2(new_n708_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n674_), .A2(new_n652_), .A3(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n786_), .A2(new_n778_), .A3(new_n636_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n784_), .A2(new_n787_), .ZN(G1332gat));
  OAI21_X1  g587(.A(G64gat), .B1(new_n786_), .B2(new_n634_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT48), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n634_), .A2(G64gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n782_), .B2(new_n791_), .ZN(G1333gat));
  OAI21_X1  g591(.A(G71gat), .B1(new_n786_), .B2(new_n663_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT49), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n663_), .A2(G71gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n782_), .B2(new_n795_), .ZN(G1334gat));
  OR3_X1    g595(.A1(new_n782_), .A2(G78gat), .A3(new_n628_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G78gat), .B1(new_n786_), .B2(new_n628_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(KEYINPUT50), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(KEYINPUT50), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(G1335gat));
  NOR2_X1   g600(.A1(new_n780_), .A2(new_n330_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n756_), .A2(new_n652_), .A3(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n803_), .A2(new_n233_), .A3(new_n636_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n651_), .A2(new_n709_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n781_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n781_), .A2(KEYINPUT115), .A3(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n641_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n233_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(KEYINPUT116), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(KEYINPUT116), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n804_), .B1(new_n813_), .B2(new_n814_), .ZN(G1336gat));
  OAI21_X1  g614(.A(G92gat), .B1(new_n803_), .B2(new_n634_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n810_), .A2(new_n234_), .A3(new_n603_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1337gat));
  NAND4_X1  g617(.A1(new_n810_), .A2(new_n435_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n819_));
  INV_X1    g618(.A(G99gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n803_), .A2(new_n663_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g622(.A1(new_n628_), .A2(G106gat), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(G106gat), .C1(new_n803_), .C2(new_n628_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n652_), .A2(new_n802_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n628_), .B(new_n829_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n830_), .B2(new_n254_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n826_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n832_), .B(new_n834_), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n213_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n216_), .A2(new_n837_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n222_), .B(new_n838_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n223_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n308_), .A2(new_n836_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n840_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT121), .B1(new_n307_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n291_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n286_), .A2(KEYINPUT55), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n289_), .A2(KEYINPUT120), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n305_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n850_), .A3(KEYINPUT56), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n848_), .B2(new_n850_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n841_), .B(new_n843_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(KEYINPUT58), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n850_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n851_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n856_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n843_), .A4(new_n841_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n857_), .A2(new_n715_), .A3(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n780_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n860_), .B2(new_n851_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n842_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n364_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT57), .B(new_n364_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n864_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n708_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n785_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT118), .B1(new_n780_), .B2(new_n708_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n715_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n879_), .A2(new_n651_), .A3(new_n880_), .A4(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n651_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n883_), .A2(new_n715_), .B1(KEYINPUT119), .B2(KEYINPUT54), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n873_), .A2(new_n885_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n635_), .A2(new_n636_), .A3(new_n663_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT123), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(G113gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n780_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n886_), .A2(KEYINPUT59), .A3(new_n888_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n228_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n896_), .B2(new_n891_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n651_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n890_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n651_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n898_), .ZN(G1341gat));
  NAND3_X1  g701(.A1(new_n890_), .A2(new_n420_), .A3(new_n330_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n708_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n420_), .ZN(G1342gat));
  NAND3_X1  g704(.A1(new_n890_), .A2(new_n418_), .A3(new_n363_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n880_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n418_), .ZN(G1343gat));
  AOI22_X1  g707(.A1(new_n872_), .A2(new_n708_), .B1(new_n884_), .B2(new_n882_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n435_), .A2(new_n628_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n636_), .A2(new_n603_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OR3_X1    g713(.A1(new_n914_), .A2(G141gat), .A3(new_n228_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G141gat), .B1(new_n914_), .B2(new_n228_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1344gat));
  OR3_X1    g716(.A1(new_n914_), .A2(G148gat), .A3(new_n651_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G148gat), .B1(new_n914_), .B2(new_n651_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n912_), .A2(new_n330_), .A3(new_n913_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1346gat));
  NOR3_X1   g722(.A1(new_n914_), .A2(new_n460_), .A3(new_n719_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n912_), .A2(new_n363_), .A3(new_n913_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n460_), .B2(new_n925_), .ZN(G1347gat));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n641_), .A2(new_n634_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n929_), .B2(new_n663_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(KEYINPUT124), .A3(new_n435_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n505_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n886_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933_), .B2(new_n228_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n933_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n937_), .A2(new_n378_), .A3(new_n380_), .A4(new_n780_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT62), .B(G169gat), .C1(new_n933_), .C2(new_n228_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(new_n938_), .A3(new_n939_), .ZN(G1348gat));
  NOR2_X1   g739(.A1(new_n933_), .A2(new_n651_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n381_), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n933_), .A2(new_n708_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(G183gat), .ZN(new_n944_));
  INV_X1    g743(.A(new_n394_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n943_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n933_), .B2(new_n880_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n363_), .A2(new_n553_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n933_), .B2(new_n948_), .ZN(G1351gat));
  NOR3_X1   g748(.A1(new_n909_), .A2(new_n911_), .A3(new_n929_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n780_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G197gat), .ZN(G1352gat));
  OAI211_X1 g751(.A(new_n950_), .B(new_n652_), .C1(KEYINPUT125), .C2(new_n476_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n950_), .A2(new_n652_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(KEYINPUT125), .B(G204gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(G1353gat));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n330_), .B1(new_n957_), .B2(new_n470_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(KEYINPUT126), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n950_), .A2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n957_), .A2(new_n470_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1354gat));
  NOR2_X1   g761(.A1(new_n364_), .A2(G218gat), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n886_), .A2(new_n910_), .A3(new_n928_), .A4(new_n963_), .ZN(new_n964_));
  NOR4_X1   g763(.A1(new_n909_), .A2(new_n880_), .A3(new_n911_), .A4(new_n929_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n965_), .B2(new_n468_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  OAI211_X1 g767(.A(KEYINPUT127), .B(new_n964_), .C1(new_n965_), .C2(new_n468_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1355gat));
endmodule


