//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n209_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT65), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  AND2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT9), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n221_), .B2(new_n215_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n205_), .B(new_n208_), .C1(new_n217_), .C2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT68), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n203_), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n225_), .B(new_n228_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n219_), .A2(new_n220_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n212_), .A2(KEYINPUT66), .A3(new_n213_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT67), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(new_n214_), .B2(new_n216_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n221_), .A2(new_n218_), .A3(new_n215_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(new_n205_), .A4(new_n208_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n228_), .A2(new_n225_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n232_), .B1(new_n204_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n235_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n224_), .A2(new_n238_), .A3(new_n243_), .A4(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G57gat), .B(G64gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT11), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G78gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n252_), .A2(KEYINPUT11), .ZN(new_n256_));
  XOR2_X1   g055(.A(G71gat), .B(G78gat), .Z(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT11), .A3(new_n252_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT12), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n259_), .ZN(new_n262_));
  AOI221_X4 g061(.A(new_n204_), .B1(new_n206_), .B2(new_n207_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n247_), .A2(new_n248_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n251_), .A2(new_n261_), .B1(new_n265_), .B2(new_n260_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n223_), .A2(new_n259_), .A3(new_n248_), .A4(new_n247_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT69), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n267_), .A2(KEYINPUT69), .A3(new_n268_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n267_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  NOR2_X1   g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT71), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n275_), .A2(new_n280_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT73), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(new_n288_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT92), .ZN(new_n296_));
  INV_X1    g095(.A(G155gat), .ZN(new_n297_));
  INV_X1    g096(.A(G162gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT92), .B1(G155gat), .B2(G162gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT93), .A4(new_n302_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G141gat), .B(G148gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT3), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT2), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT94), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n299_), .A2(new_n302_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT94), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n316_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n323_), .A2(new_n300_), .A3(new_n325_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n310_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G120gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(G127gat), .A2(G134gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G127gat), .A2(G134gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT90), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G127gat), .ZN(new_n334_));
  INV_X1    g133(.A(G134gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT90), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G127gat), .A2(G134gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G113gat), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n333_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n333_), .B2(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n330_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT90), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n337_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n345_));
  OAI21_X1  g144(.A(G113gat), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n333_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(G120gat), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n329_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n310_), .A2(new_n328_), .A3(new_n348_), .A4(new_n343_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT4), .A4(new_n352_), .ZN(new_n353_));
  AND4_X1   g152(.A1(new_n310_), .A2(new_n328_), .A3(new_n348_), .A4(new_n343_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n310_), .A2(new_n328_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT98), .B1(new_n350_), .B2(KEYINPUT4), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT100), .ZN(new_n363_));
  NOR4_X1   g162(.A1(new_n354_), .A2(new_n355_), .A3(new_n363_), .A4(new_n361_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n354_), .A2(new_n355_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT100), .B1(new_n372_), .B2(new_n360_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n362_), .A2(new_n365_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G64gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(G64gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n211_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G92gat), .A3(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(KEYINPUT88), .A2(G169gat), .A3(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393_));
  INV_X1    g192(.A(G169gat), .ZN(new_n394_));
  INV_X1    g193(.A(G176gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT87), .B1(G169gat), .B2(G176gat), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n392_), .A2(KEYINPUT24), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n399_));
  AND2_X1   g198(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n402_));
  OAI22_X1  g201(.A1(new_n399_), .A2(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404_));
  INV_X1    g203(.A(new_n397_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(KEYINPUT87), .A2(G169gat), .A3(G176gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n398_), .A2(new_n403_), .A3(new_n407_), .A4(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n414_), .A3(new_n411_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT22), .B(G169gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n395_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n410_), .A2(new_n414_), .A3(KEYINPUT89), .A4(new_n411_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n417_), .A2(new_n392_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G211gat), .B(G218gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G197gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(G204gat), .ZN(new_n425_));
  INV_X1    g224(.A(G204gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(G197gat), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n423_), .B(KEYINPUT21), .C1(new_n425_), .C2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G197gat), .B(G204gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT21), .B1(new_n425_), .B2(new_n427_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n422_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n413_), .A2(new_n421_), .A3(new_n428_), .A4(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n396_), .A2(KEYINPUT24), .A3(new_n397_), .A4(new_n388_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n407_), .A2(new_n435_), .A3(new_n412_), .A4(new_n403_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n419_), .A2(new_n392_), .A3(new_n415_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n428_), .A2(new_n433_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G226gat), .A2(G233gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT19), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n434_), .A2(new_n440_), .A3(KEYINPUT20), .A4(new_n442_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n413_), .A2(new_n421_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n438_), .A2(new_n439_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n387_), .B(new_n443_), .C1(new_n447_), .C2(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT97), .ZN(new_n449_));
  INV_X1    g248(.A(new_n387_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n444_), .A2(new_n446_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n445_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n442_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n442_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n413_), .A2(new_n421_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n439_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT20), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n456_), .B1(new_n459_), .B2(new_n445_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT97), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n387_), .A4(new_n443_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n449_), .A2(new_n455_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n372_), .A2(new_n361_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n371_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n373_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n376_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(new_n371_), .A3(new_n365_), .A4(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n377_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n450_), .A2(KEYINPUT32), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n447_), .A2(new_n456_), .ZN(new_n473_));
  AND4_X1   g272(.A1(KEYINPUT20), .A2(new_n434_), .A3(new_n440_), .A4(new_n456_), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT32), .B(new_n450_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n371_), .B1(new_n467_), .B2(new_n365_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n350_), .A2(KEYINPUT4), .A3(new_n352_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n351_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n360_), .B1(new_n479_), .B2(new_n353_), .ZN(new_n480_));
  NOR4_X1   g279(.A1(new_n480_), .A2(new_n370_), .A3(new_n364_), .A4(new_n373_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n472_), .B(new_n475_), .C1(new_n476_), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n470_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G22gat), .B(G50gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n327_), .A2(new_n300_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n324_), .B1(new_n322_), .B2(KEYINPUT94), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n488_), .A2(new_n489_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT29), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n487_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  AND4_X1   g291(.A1(new_n491_), .A2(new_n310_), .A3(new_n328_), .A4(new_n487_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n485_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n486_), .B1(new_n329_), .B2(KEYINPUT29), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n484_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G78gat), .B(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n329_), .A2(KEYINPUT29), .B1(new_n428_), .B2(new_n433_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G228gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n500_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n494_), .A2(new_n497_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G71gat), .B(G99gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT30), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G227gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G15gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n512_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G43gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n413_), .A2(new_n517_), .A3(new_n421_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n413_), .B2(new_n421_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n516_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(KEYINPUT91), .A3(new_n523_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n349_), .B(KEYINPUT31), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n510_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n483_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n476_), .A2(new_n481_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n387_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n535_), .A2(KEYINPUT27), .A3(new_n455_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n463_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n508_), .A2(new_n531_), .A3(new_n509_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n530_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n509_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n541_), .B2(new_n507_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n534_), .B(new_n538_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n533_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n295_), .A2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G15gat), .B(G22gat), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(KEYINPUT80), .A2(G8gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(KEYINPUT80), .A2(G8gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(G1gat), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT81), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT14), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n550_), .B2(KEYINPUT14), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n547_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G1gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(KEYINPUT14), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT81), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n546_), .B1(new_n558_), .B2(new_n552_), .ZN(new_n559_));
  INV_X1    g358(.A(G1gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n561_), .A3(G8gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(G8gat), .B1(new_n556_), .B2(new_n561_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT82), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n259_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n565_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G183gat), .ZN(new_n573_));
  INV_X1    g372(.A(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  OR4_X1    g374(.A1(KEYINPUT83), .A2(new_n569_), .A3(new_n570_), .A4(new_n575_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n569_), .A2(KEYINPUT83), .B1(new_n570_), .B2(new_n575_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(G29gat), .A2(G36gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G29gat), .A2(G36gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n517_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G43gat), .B1(new_n585_), .B2(new_n581_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n584_), .A2(new_n586_), .A3(G50gat), .ZN(new_n587_));
  AOI21_X1  g386(.A(G50gat), .B1(new_n584_), .B2(new_n586_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT15), .ZN(new_n590_));
  AND4_X1   g389(.A1(new_n248_), .A2(new_n223_), .A3(new_n589_), .A4(new_n247_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n251_), .A2(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT74), .Z(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT34), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n223_), .A2(new_n248_), .A3(new_n247_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n589_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT75), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n593_), .A2(new_n597_), .A3(new_n600_), .A4(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G134gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n298_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT77), .Z(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT76), .B(new_n597_), .C1(new_n593_), .C2(new_n600_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT76), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n251_), .A2(new_n590_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n591_), .A2(new_n592_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n600_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n597_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n603_), .B(new_n609_), .C1(new_n610_), .C2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n618_));
  INV_X1    g417(.A(new_n603_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT76), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n614_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n606_), .B(KEYINPUT36), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n617_), .B(new_n618_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(KEYINPUT78), .A3(new_n609_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT37), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT79), .B(KEYINPUT37), .Z(new_n629_));
  OAI211_X1 g428(.A(new_n617_), .B(new_n629_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT86), .ZN(new_n632_));
  INV_X1    g431(.A(G8gat), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n555_), .A2(G1gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n559_), .A2(new_n560_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n599_), .B1(new_n636_), .B2(new_n562_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT84), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT85), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n589_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT85), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT84), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n565_), .A2(new_n599_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n639_), .A2(new_n642_), .A3(new_n565_), .A4(new_n599_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n565_), .A2(new_n590_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n646_), .A3(new_n640_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(new_n394_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(new_n424_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n649_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n632_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n649_), .A2(new_n651_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n654_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n649_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(KEYINPUT86), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n545_), .A2(new_n580_), .A3(new_n631_), .A4(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT102), .Z(new_n666_));
  INV_X1    g465(.A(new_n534_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n560_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT38), .ZN(new_n669_));
  INV_X1    g468(.A(new_n295_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n656_), .A2(new_n657_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n617_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n533_), .B2(new_n543_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT103), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n580_), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n677_), .B2(new_n534_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  OAI221_X1 g480(.A(G8gat), .B1(new_n680_), .B2(new_n681_), .C1(new_n677_), .C2(new_n538_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n548_), .A2(new_n549_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n538_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n666_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n677_), .B2(new_n540_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT41), .Z(new_n692_));
  INV_X1    g491(.A(G15gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n666_), .A2(new_n693_), .A3(new_n531_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1326gat));
  INV_X1    g494(.A(G22gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n666_), .A2(new_n696_), .A3(new_n510_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n510_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G22gat), .B1(new_n677_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n580_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n674_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n295_), .A2(new_n544_), .A3(new_n664_), .A4(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n667_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n628_), .A2(new_n630_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n544_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n544_), .A2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT43), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n544_), .A2(new_n709_), .A3(KEYINPUT105), .A4(new_n708_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n671_), .ZN(new_n717_));
  AND4_X1   g516(.A1(new_n702_), .A2(new_n292_), .A3(new_n717_), .A4(new_n294_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n719_), .A2(G29gat), .A3(new_n667_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n718_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n707_), .B1(new_n720_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n705_), .A2(G36gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n686_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(KEYINPUT45), .A3(new_n686_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n716_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT44), .B1(new_n716_), .B2(new_n718_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n538_), .ZN(new_n735_));
  INV_X1    g534(.A(G36gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT106), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n723_), .A2(new_n686_), .A3(new_n719_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n739_), .A3(G36gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n732_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n725_), .B(new_n726_), .C1(new_n741_), .C2(KEYINPUT107), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT46), .B1(new_n741_), .B2(new_n725_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n732_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n538_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n745_));
  AOI211_X1 g544(.A(KEYINPUT106), .B(new_n736_), .C1(new_n745_), .C2(new_n719_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n739_), .B1(new_n738_), .B2(G36gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT108), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n742_), .B1(new_n743_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(G1329gat));
  AOI21_X1  g551(.A(G43gat), .B1(new_n706_), .B2(new_n531_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n733_), .A2(new_n734_), .A3(new_n517_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n531_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g555(.A(G50gat), .B1(new_n706_), .B2(new_n510_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n723_), .A2(G50gat), .A3(new_n719_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n510_), .ZN(G1331gat));
  NOR2_X1   g558(.A1(new_n295_), .A2(new_n717_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n544_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(new_n702_), .A3(new_n709_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n667_), .ZN(new_n763_));
  AND4_X1   g562(.A1(new_n580_), .A2(new_n676_), .A3(new_n670_), .A4(new_n663_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n667_), .A2(G57gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n764_), .B2(new_n765_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n764_), .B2(new_n686_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT48), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n762_), .A2(new_n767_), .A3(new_n686_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n764_), .B2(new_n531_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT49), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n772_), .A3(new_n531_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  INV_X1    g575(.A(G78gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n764_), .B2(new_n510_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT50), .Z(new_n779_));
  NAND2_X1  g578(.A1(new_n510_), .A2(new_n777_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT109), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n762_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n761_), .A2(new_n703_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n667_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n760_), .A2(new_n702_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT110), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n716_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n534_), .A2(new_n210_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(G1336gat));
  AOI21_X1  g590(.A(G92gat), .B1(new_n784_), .B2(new_n686_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n538_), .A2(new_n211_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n789_), .B2(new_n793_), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n788_), .B2(new_n540_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n784_), .A2(new_n206_), .A3(new_n531_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g597(.A1(new_n784_), .A2(new_n207_), .A3(new_n510_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n510_), .A3(new_n716_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(G106gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT53), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n799_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n266_), .A2(new_n811_), .A3(new_n267_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n273_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n251_), .A2(new_n261_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n265_), .A2(new_n260_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n270_), .A2(new_n269_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n817_), .A2(new_n818_), .B1(KEYINPUT111), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT111), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n271_), .A2(KEYINPUT111), .A3(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n814_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n280_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(new_n280_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n284_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n275_), .A2(new_n283_), .A3(new_n280_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n826_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n650_), .A2(new_n640_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n650_), .A2(KEYINPUT113), .A3(new_n640_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n647_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n654_), .A3(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n661_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n831_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n810_), .B1(new_n840_), .B2(new_n631_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n824_), .A2(new_n280_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT56), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n824_), .A2(new_n825_), .A3(new_n280_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n285_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n661_), .A2(new_n838_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT58), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT115), .B(new_n709_), .C1(new_n847_), .C2(KEYINPUT58), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n841_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n671_), .A2(new_n845_), .B1(new_n289_), .B2(new_n846_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT116), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n673_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n855_), .B2(new_n852_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n851_), .A2(new_n673_), .A3(new_n856_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n850_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n702_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n663_), .A2(new_n580_), .A3(new_n291_), .A4(new_n631_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT59), .B1(new_n866_), .B2(KEYINPUT118), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n667_), .A2(new_n538_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n542_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n864_), .B1(new_n860_), .B2(new_n702_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n542_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n868_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n877_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n340_), .B(new_n663_), .C1(new_n871_), .C2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n872_), .A2(new_n873_), .A3(new_n671_), .A4(new_n868_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(G113gat), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT117), .B(new_n340_), .C1(new_n870_), .C2(new_n671_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n809_), .B1(new_n879_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n871_), .A2(new_n878_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(G113gat), .A3(new_n664_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n887_), .A2(KEYINPUT119), .A3(new_n883_), .A4(new_n882_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1340gat));
  AND2_X1   g688(.A1(new_n330_), .A2(KEYINPUT60), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT60), .B1(new_n670_), .B2(new_n330_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n870_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n295_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n330_), .ZN(G1341gat));
  AOI21_X1  g695(.A(G127gat), .B1(new_n874_), .B2(new_n580_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n702_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g698(.A(G134gat), .B1(new_n874_), .B2(new_n674_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n631_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(G134gat), .ZN(G1343gat));
  NOR4_X1   g701(.A1(new_n872_), .A2(new_n531_), .A3(new_n698_), .A4(new_n868_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n717_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n670_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT121), .B(G148gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n903_), .A2(new_n580_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  AOI21_X1  g710(.A(G162gat), .B1(new_n903_), .B2(new_n674_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n631_), .A2(new_n298_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n913_), .ZN(G1347gat));
  NOR3_X1   g713(.A1(new_n872_), .A2(new_n667_), .A3(new_n873_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n915_), .A2(new_n686_), .A3(new_n717_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n916_), .A2(new_n917_), .A3(G169gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n916_), .B2(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n686_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n717_), .A2(new_n418_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(KEYINPUT122), .Z(new_n922_));
  OAI22_X1  g721(.A1(new_n918_), .A2(new_n919_), .B1(new_n920_), .B2(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n920_), .A2(new_n295_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n395_), .ZN(G1349gat));
  NOR2_X1   g724(.A1(new_n920_), .A2(new_n702_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n927_));
  INV_X1    g726(.A(G183gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(new_n926_), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n915_), .A2(new_n686_), .A3(new_n709_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n930_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT123), .B1(new_n930_), .B2(G190gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n674_), .B1(new_n402_), .B2(new_n401_), .ZN(new_n933_));
  OAI22_X1  g732(.A1(new_n931_), .A2(new_n932_), .B1(new_n920_), .B2(new_n933_), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n539_), .A2(new_n534_), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT124), .Z(new_n936_));
  NAND3_X1  g735(.A1(new_n866_), .A2(new_n686_), .A3(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT125), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n938_), .A2(G197gat), .A3(new_n717_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G197gat), .B1(new_n938_), .B2(new_n717_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n670_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(G204gat), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n938_), .A2(new_n426_), .A3(new_n670_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1353gat));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n574_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n580_), .B1(new_n947_), .B2(new_n574_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT126), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n938_), .A2(new_n948_), .A3(new_n950_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n948_), .B1(new_n938_), .B2(new_n950_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n938_), .B2(new_n674_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n938_), .A2(new_n709_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(G218gat), .B2(new_n956_), .ZN(G1355gat));
endmodule


