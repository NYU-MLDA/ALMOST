//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n841_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT31), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT79), .B1(new_n208_), .B2(KEYINPUT26), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n207_), .B(new_n209_), .C1(new_n210_), .C2(KEYINPUT79), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n211_), .A2(new_n213_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n222_), .B(new_n223_), .C1(G183gat), .C2(G190gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n225_));
  OR3_X1    g024(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(G15gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT30), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n235_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n206_), .B1(new_n239_), .B2(KEYINPUT80), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(KEYINPUT80), .B2(new_n239_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n242_), .A3(new_n206_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G78gat), .B(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G197gat), .ZN(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G204gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT85), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n250_), .B(KEYINPUT87), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n248_), .B(KEYINPUT86), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n252_), .B(new_n253_), .C1(KEYINPUT21), .C2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n253_), .A2(new_n246_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G228gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n270_));
  OR2_X1    g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n268_), .A2(new_n267_), .A3(KEYINPUT1), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n265_), .B(new_n266_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n265_), .B(KEYINPUT2), .ZN(new_n278_));
  OR4_X1    g077(.A1(KEYINPUT82), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT3), .B1(new_n266_), .B2(KEYINPUT82), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n277_), .B1(KEYINPUT83), .B2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(KEYINPUT83), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n274_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n264_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n260_), .A2(KEYINPUT89), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n257_), .A2(new_n288_), .A3(new_n259_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n262_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n245_), .B1(new_n286_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n289_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n288_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n297_), .A2(new_n263_), .B1(new_n264_), .B2(new_n285_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n245_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n301_));
  XOR2_X1   g100(.A(G22gat), .B(G50gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT28), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n301_), .B(new_n303_), .ZN(new_n304_));
  AND4_X1   g103(.A1(KEYINPUT90), .A2(new_n294_), .A3(new_n300_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT90), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n306_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n307_), .A2(new_n304_), .B1(new_n294_), .B2(new_n300_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n257_), .A2(new_n259_), .A3(new_n227_), .A4(new_n220_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n227_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n210_), .A2(new_n207_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n312_), .A2(new_n218_), .A3(new_n213_), .A4(new_n219_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT92), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n314_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n311_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(KEYINPUT20), .B(new_n310_), .C1(new_n261_), .C2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n261_), .A2(new_n317_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n260_), .A2(new_n228_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n324_), .A2(KEYINPUT20), .A3(new_n321_), .A4(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G64gat), .B(G92gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n323_), .A2(new_n331_), .A3(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n284_), .A2(new_n204_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n337_));
  INV_X1    g136(.A(new_n204_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n274_), .C1(new_n283_), .C2(new_n282_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n284_), .A2(new_n337_), .A3(new_n204_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G1gat), .B(G29gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n342_), .A2(KEYINPUT4), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n284_), .A2(new_n204_), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n343_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT98), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n352_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n353_), .A2(KEYINPUT98), .A3(new_n343_), .A4(new_n355_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n335_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n342_), .A2(new_n343_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n355_), .A2(new_n344_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n361_), .B(new_n350_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT33), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT96), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n344_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n364_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n353_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT33), .A4(new_n350_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n365_), .A2(new_n374_), .A3(new_n366_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n360_), .B(new_n373_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n318_), .A2(new_n322_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT100), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n313_), .A2(new_n227_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT99), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n295_), .A2(new_n296_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n379_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n290_), .C2(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n325_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n378_), .B1(new_n386_), .B2(new_n322_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT101), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT101), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n381_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n392_), .A2(new_n379_), .B1(new_n260_), .B2(new_n228_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n321_), .B1(new_n393_), .B2(new_n385_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n390_), .B(new_n391_), .C1(new_n394_), .C2(new_n378_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n327_), .A2(new_n391_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n363_), .A2(new_n364_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n351_), .B1(new_n397_), .B2(new_n368_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n398_), .B2(new_n365_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n389_), .A2(new_n395_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n309_), .B1(new_n377_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  INV_X1    g201(.A(new_n334_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n331_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT102), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n335_), .A2(KEYINPUT102), .A3(new_n402_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT27), .B(new_n334_), .C1(new_n387_), .C2(new_n331_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n398_), .A2(new_n365_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AND4_X1   g211(.A1(new_n309_), .A2(new_n409_), .A3(new_n410_), .A4(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n244_), .B1(new_n401_), .B2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n409_), .A2(new_n410_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n309_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n244_), .A2(new_n411_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G230gat), .A2(G233gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n421_), .A2(KEYINPUT9), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G99gat), .A2(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT6), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G99gat), .A3(G106gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n428_));
  INV_X1    g227(.A(G106gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G85gat), .ZN(new_n432_));
  INV_X1    g231(.A(G92gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(KEYINPUT9), .A3(new_n421_), .ZN(new_n435_));
  AND4_X1   g234(.A1(new_n422_), .A2(new_n427_), .A3(new_n431_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n421_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n429_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT8), .B(new_n438_), .C1(new_n443_), .C2(new_n427_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n427_), .A2(new_n442_), .A3(new_n441_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n438_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n437_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n424_), .A2(new_n426_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n441_), .A2(new_n442_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n447_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT8), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT64), .A3(new_n437_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n461_));
  XOR2_X1   g260(.A(G71gat), .B(G78gat), .Z(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n451_), .A2(new_n458_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n449_), .A2(new_n467_), .A3(KEYINPUT12), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n465_), .B1(new_n451_), .B2(new_n458_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT64), .B1(new_n457_), .B2(new_n437_), .ZN(new_n475_));
  AOI211_X1 g274(.A(new_n450_), .B(new_n436_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n467_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n473_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT67), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n420_), .B(new_n470_), .C1(new_n474_), .C2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(KEYINPUT65), .A3(new_n466_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n420_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n481_), .B(new_n482_), .C1(KEYINPUT65), .C2(new_n477_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT68), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT69), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT68), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n480_), .A2(new_n487_), .A3(new_n483_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G120gat), .B(G148gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT5), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G176gat), .B(G204gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  NAND4_X1  g291(.A1(new_n485_), .A2(new_n486_), .A3(new_n488_), .A4(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n480_), .A2(new_n487_), .A3(new_n483_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n487_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n492_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n480_), .A2(new_n483_), .A3(new_n496_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT69), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n493_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT13), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT13), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n493_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505_));
  INV_X1    g304(.A(G1gat), .ZN(new_n506_));
  INV_X1    g305(.A(G8gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT74), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G8gat), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G29gat), .B(G36gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT77), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n515_), .A2(new_n518_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n515_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n518_), .B(KEYINPUT15), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n520_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n528_), .B2(new_n522_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G113gat), .B(G141gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT78), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n524_), .B(new_n535_), .C1(new_n528_), .C2(new_n522_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n504_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n419_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  XOR2_X1   g340(.A(G190gat), .B(G218gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT70), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT36), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n451_), .A2(new_n458_), .A3(new_n518_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n526_), .B2(new_n449_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n547_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n546_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n554_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT71), .Z(new_n559_));
  AOI22_X1  g358(.A1(new_n555_), .A2(new_n556_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n555_), .A2(new_n556_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n541_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n559_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n565_), .A2(new_n555_), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n562_), .A2(new_n563_), .B1(new_n541_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n465_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT75), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(new_n525_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n571_), .B(new_n515_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n568_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT76), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n540_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n506_), .A3(new_n411_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT38), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n539_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n583_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n566_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n412_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n590_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n596_), .A3(new_n597_), .ZN(G1324gat));
  INV_X1    g397(.A(new_n415_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n507_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  INV_X1    g400(.A(new_n595_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n599_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n603_), .B2(G8gat), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT39), .B(new_n507_), .C1(new_n602_), .C2(new_n599_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g406(.A(new_n244_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n233_), .B1(new_n602_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(KEYINPUT41), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(new_n611_), .B2(new_n612_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n587_), .A2(G15gat), .A3(new_n244_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(G1326gat));
  OR3_X1    g415(.A1(new_n587_), .A2(G22gat), .A3(new_n416_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n602_), .A2(new_n309_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT42), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n618_), .A2(new_n619_), .A3(G22gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n618_), .B2(G22gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT104), .ZN(G1327gat));
  NOR2_X1   g422(.A1(new_n592_), .A2(new_n584_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  INV_X1    g424(.A(new_n568_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n625_), .B1(new_n419_), .B2(new_n626_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT43), .B(new_n568_), .C1(new_n414_), .C2(new_n418_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT44), .B(new_n624_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n412_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n566_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n584_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n540_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n412_), .A2(G29gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT105), .Z(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n637_), .B2(new_n639_), .ZN(G1328gat));
  NOR3_X1   g439(.A1(new_n637_), .A2(G36gat), .A3(new_n415_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n631_), .A2(new_n599_), .A3(new_n632_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(KEYINPUT106), .ZN(new_n645_));
  OAI21_X1  g444(.A(G36gat), .B1(new_n644_), .B2(KEYINPUT106), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI221_X1 g448(.A(new_n643_), .B1(KEYINPUT108), .B2(KEYINPUT46), .C1(new_n645_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  OAI21_X1  g450(.A(G43gat), .B1(new_n633_), .B2(new_n244_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n244_), .A2(G43gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n637_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1330gat));
  INV_X1    g455(.A(G50gat), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n633_), .A2(new_n657_), .A3(new_n416_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n540_), .A2(new_n309_), .A3(new_n636_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n657_), .B2(new_n659_), .ZN(G1331gat));
  AND3_X1   g459(.A1(new_n419_), .A2(new_n538_), .A3(new_n504_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n586_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n411_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n504_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n578_), .A2(new_n582_), .A3(new_n536_), .A4(new_n534_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n594_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G57gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n411_), .B2(KEYINPUT110), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(KEYINPUT110), .B2(new_n670_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n664_), .B1(new_n669_), .B2(new_n672_), .ZN(G1332gat));
  OAI21_X1  g472(.A(G64gat), .B1(new_n668_), .B2(new_n415_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT48), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n415_), .A2(G64gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n662_), .B2(new_n676_), .ZN(G1333gat));
  OAI21_X1  g476(.A(G71gat), .B1(new_n668_), .B2(new_n244_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT49), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n244_), .A2(G71gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n662_), .B2(new_n680_), .ZN(G1334gat));
  OR3_X1    g480(.A1(new_n662_), .A2(G78gat), .A3(new_n416_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n669_), .A2(new_n309_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(G78gat), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G78gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT112), .Z(G1335gat));
  NOR3_X1   g487(.A1(new_n665_), .A2(new_n584_), .A3(new_n537_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n627_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n419_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G85gat), .B1(new_n694_), .B2(new_n412_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n661_), .A2(new_n636_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT113), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n411_), .A2(new_n432_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(G1336gat));
  OAI21_X1  g500(.A(G92gat), .B1(new_n694_), .B2(new_n415_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n599_), .A2(new_n433_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n699_), .B2(new_n703_), .ZN(G1337gat));
  INV_X1    g503(.A(KEYINPUT115), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n608_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n698_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n693_), .A2(new_n608_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n708_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT114), .B1(new_n708_), .B2(G99gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n707_), .B(new_n712_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1338gat));
  OAI211_X1 g515(.A(new_n309_), .B(new_n689_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT117), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G106gat), .B1(new_n717_), .B2(new_n718_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT52), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n693_), .A2(KEYINPUT117), .A3(new_n309_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .A4(new_n719_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n698_), .A2(new_n429_), .A3(new_n309_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n726_), .A2(new_n730_), .A3(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1339gat));
  INV_X1    g531(.A(KEYINPUT59), .ZN(new_n733_));
  NOR4_X1   g532(.A1(new_n599_), .A2(new_n309_), .A3(new_n412_), .A4(new_n244_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n735_), .B2(KEYINPUT124), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(KEYINPUT124), .B2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n528_), .A2(new_n522_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n520_), .A2(new_n523_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n533_), .B1(new_n739_), .B2(new_n521_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n529_), .A2(new_n533_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n498_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n472_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n477_), .A2(KEYINPUT67), .A3(new_n478_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n470_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT120), .A3(new_n482_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT120), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n469_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n420_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n480_), .A2(KEYINPUT55), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n749_), .A2(new_n753_), .A3(new_n420_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n751_), .A2(new_n755_), .A3(KEYINPUT121), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT121), .B1(new_n751_), .B2(new_n755_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n492_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT56), .B(new_n492_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n742_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n626_), .B1(new_n762_), .B2(KEYINPUT58), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n764_), .B(new_n742_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n493_), .B(new_n741_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT123), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n537_), .A2(new_n498_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT122), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT122), .B(new_n769_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n635_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n766_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT57), .B(new_n635_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n584_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n666_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n779_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n781_), .A2(new_n782_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n779_), .A3(new_n784_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT119), .B(KEYINPUT54), .C1(new_n781_), .C2(new_n782_), .ZN(new_n790_));
  OAI22_X1  g589(.A1(new_n785_), .A2(new_n790_), .B1(new_n782_), .B2(new_n781_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n737_), .B1(new_n778_), .B2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n763_), .A2(new_n765_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT123), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n767_), .B(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n769_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT120), .B1(new_n746_), .B2(new_n482_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n749_), .A2(new_n748_), .A3(new_n420_), .ZN(new_n799_));
  AND4_X1   g598(.A1(new_n753_), .A2(new_n745_), .A3(new_n420_), .A4(new_n470_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n753_), .B1(new_n749_), .B2(new_n420_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n798_), .A2(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT121), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n751_), .A2(new_n755_), .A3(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n492_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n759_), .B(new_n496_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n797_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n796_), .B1(new_n809_), .B2(KEYINPUT122), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n770_), .A2(new_n771_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n566_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n794_), .B1(new_n812_), .B2(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(new_n777_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n583_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n792_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n735_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n537_), .B(new_n793_), .C1(new_n817_), .C2(new_n733_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G113gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n734_), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n821_), .A2(G113gat), .A3(new_n538_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n822_), .ZN(G1340gat));
  OAI211_X1 g622(.A(new_n504_), .B(new_n793_), .C1(new_n817_), .C2(new_n733_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G120gat), .ZN(new_n825_));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n665_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n817_), .B(new_n827_), .C1(KEYINPUT60), .C2(new_n826_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1341gat));
  OAI211_X1 g628(.A(new_n584_), .B(new_n793_), .C1(new_n817_), .C2(new_n733_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G127gat), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n821_), .A2(G127gat), .A3(new_n583_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1342gat));
  OAI211_X1 g632(.A(new_n626_), .B(new_n793_), .C1(new_n817_), .C2(new_n733_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G134gat), .ZN(new_n835_));
  OR3_X1    g634(.A1(new_n821_), .A2(G134gat), .A3(new_n635_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1343gat));
  NOR4_X1   g636(.A1(new_n599_), .A2(new_n416_), .A3(new_n412_), .A4(new_n608_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n820_), .A2(new_n537_), .A3(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g639(.A1(new_n820_), .A2(new_n504_), .A3(new_n838_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g641(.A1(new_n820_), .A2(new_n584_), .A3(new_n838_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT61), .B(G155gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1346gat));
  AND4_X1   g644(.A1(G162gat), .A2(new_n820_), .A3(new_n626_), .A4(new_n838_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n566_), .B(new_n838_), .C1(new_n778_), .C2(new_n792_), .ZN(new_n847_));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT125), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT125), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n846_), .B1(new_n850_), .B2(new_n852_), .ZN(G1347gat));
  NAND3_X1  g652(.A1(new_n599_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT126), .B1(new_n820_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n774_), .A2(new_n775_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n777_), .A3(new_n794_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n792_), .B1(new_n858_), .B2(new_n583_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n854_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT22), .B(G169gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n537_), .A2(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n537_), .B(new_n855_), .C1(new_n778_), .C2(new_n792_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n865_), .A2(new_n866_), .A3(G169gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n865_), .B2(G169gat), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n862_), .A2(new_n864_), .B1(new_n867_), .B2(new_n868_), .ZN(G1348gat));
  NAND2_X1  g668(.A1(new_n504_), .A2(new_n217_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n859_), .A2(new_n665_), .A3(new_n854_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n862_), .A2(new_n870_), .B1(new_n217_), .B2(new_n871_), .ZN(G1349gat));
  OAI21_X1  g671(.A(new_n860_), .B1(new_n859_), .B2(new_n854_), .ZN(new_n873_));
  OAI211_X1 g672(.A(KEYINPUT126), .B(new_n855_), .C1(new_n778_), .C2(new_n792_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n583_), .A2(new_n207_), .ZN(new_n876_));
  INV_X1    g675(.A(G183gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n820_), .A2(new_n584_), .A3(new_n855_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n875_), .A2(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1350gat));
  AND2_X1   g678(.A1(new_n566_), .A2(new_n210_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n568_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n208_), .B2(new_n882_), .ZN(G1351gat));
  XOR2_X1   g682(.A(KEYINPUT127), .B(G197gat), .Z(new_n884_));
  NOR4_X1   g683(.A1(new_n415_), .A2(new_n416_), .A3(new_n411_), .A4(new_n608_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n820_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(new_n538_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n249_), .A2(KEYINPUT127), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n820_), .A2(new_n537_), .A3(new_n885_), .A4(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1352gat));
  NAND3_X1  g689(.A1(new_n820_), .A2(new_n504_), .A3(new_n885_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g691(.A(KEYINPUT63), .B(G211gat), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n820_), .A2(new_n584_), .A3(new_n885_), .A4(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n886_), .A2(new_n583_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(G1354gat));
  OAI21_X1  g696(.A(G218gat), .B1(new_n886_), .B2(new_n568_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n635_), .A2(G218gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n886_), .B2(new_n899_), .ZN(G1355gat));
endmodule


