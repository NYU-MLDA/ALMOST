//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT67), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n206_), .B(new_n208_), .C1(new_n209_), .C2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT65), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT65), .B1(new_n214_), .B2(new_n216_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n214_), .A2(new_n216_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  INV_X1    g021(.A(G99gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n205_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n207_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT8), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  INV_X1    g028(.A(new_n225_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G85gat), .B(G92gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT8), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n228_), .A2(new_n229_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n227_), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n220_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n242_));
  XOR2_X1   g041(.A(G71gat), .B(G78gat), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n203_), .B1(new_n238_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G230gat), .A2(G233gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n214_), .A2(new_n216_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n234_), .B1(new_n232_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT8), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n229_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n233_), .A2(new_n235_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n237_), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n212_), .A2(new_n219_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n246_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n256_), .A2(new_n257_), .B1(KEYINPUT67), .B2(new_n202_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n202_), .A2(KEYINPUT67), .ZN(new_n259_));
  AOI211_X1 g058(.A(new_n259_), .B(new_n246_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n247_), .B(new_n248_), .C1(new_n258_), .C2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n238_), .A2(new_n246_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n257_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n248_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G120gat), .B(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G176gat), .B(G204gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT13), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT68), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G232gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT34), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G29gat), .B(G36gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT70), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT71), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G43gat), .B(G50gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n286_), .A2(KEYINPUT70), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(KEYINPUT70), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n289_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n289_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n291_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n238_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n283_), .A2(new_n284_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT15), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n296_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n289_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n298_), .A2(KEYINPUT15), .A3(new_n294_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n238_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n285_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n303_), .A2(new_n304_), .A3(new_n302_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT15), .B1(new_n298_), .B2(new_n294_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n256_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n285_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n300_), .A4(new_n299_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G190gat), .B(G218gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT72), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G134gat), .B(G162gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT36), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n308_), .A2(new_n313_), .A3(KEYINPUT73), .A4(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n317_), .B(new_n318_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT37), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n329_), .B(new_n326_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G1gat), .ZN(new_n332_));
  INV_X1    g131(.A(G8gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT14), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n334_), .A2(KEYINPUT74), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(KEYINPUT74), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G15gat), .B(G22gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G1gat), .B(G8gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n335_), .A2(new_n341_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(new_n246_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G231gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G127gat), .B(G155gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT17), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n351_), .B(KEYINPUT17), .Z(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n346_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n331_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n280_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT19), .ZN(new_n363_));
  XOR2_X1   g162(.A(G211gat), .B(G218gat), .Z(new_n364_));
  INV_X1    g163(.A(G197gat), .ZN(new_n365_));
  INV_X1    g164(.A(G204gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT82), .B(G197gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n366_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT21), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n365_), .B2(G204gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n368_), .B2(G204gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n375_), .A2(G197gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n365_), .A2(KEYINPUT82), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n372_), .B(new_n366_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n378_), .A3(KEYINPUT21), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n371_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n369_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT84), .B(new_n367_), .C1(new_n368_), .C2(new_n366_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n364_), .A2(KEYINPUT21), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G169gat), .ZN(new_n387_));
  INV_X1    g186(.A(G176gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT78), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT23), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n394_), .B(new_n395_), .C1(G183gat), .C2(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n387_), .A2(new_n397_), .A3(new_n388_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n390_), .A2(new_n391_), .A3(new_n396_), .A4(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT25), .B(G183gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n401_));
  INV_X1    g200(.A(G190gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(KEYINPUT26), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT26), .B(G190gat), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n400_), .B(new_n403_), .C1(new_n404_), .C2(new_n401_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n392_), .B(KEYINPUT23), .ZN(new_n406_));
  NOR3_X1   g205(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n409_), .B2(new_n391_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n399_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n386_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n391_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT88), .B(new_n391_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n400_), .A2(new_n404_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n416_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n414_), .A3(new_n421_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n406_), .A2(KEYINPUT89), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT89), .B1(new_n406_), .B2(new_n426_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n423_), .B(new_n424_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n389_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n429_), .A2(new_n430_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n363_), .B1(new_n413_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n386_), .B2(new_n412_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n363_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n429_), .A2(new_n380_), .A3(new_n385_), .A4(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(KEYINPUT90), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n434_), .A2(new_n439_), .A3(new_n435_), .A4(new_n436_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n361_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  INV_X1    g241(.A(new_n361_), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n413_), .A2(new_n431_), .A3(new_n363_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n436_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n363_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n441_), .A2(new_n442_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n438_), .A2(new_n361_), .A3(new_n440_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n441_), .B2(KEYINPUT91), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n438_), .A2(new_n440_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n451_), .A2(KEYINPUT91), .A3(new_n443_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT100), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(KEYINPUT100), .B(new_n442_), .C1(new_n450_), .C2(new_n452_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n448_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G113gat), .B(G120gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G134gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G127gat), .ZN(new_n462_));
  INV_X1    g261(.A(G127gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G134gat), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n462_), .A2(new_n464_), .A3(KEYINPUT79), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT79), .B1(new_n462_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n460_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n463_), .A2(G134gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n461_), .A2(G127gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n464_), .A3(KEYINPUT79), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n459_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G141gat), .A2(G148gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT3), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n479_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n477_), .B1(KEYINPUT1), .B2(new_n475_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n475_), .A2(KEYINPUT1), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G141gat), .B(G148gat), .Z(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n474_), .B1(new_n490_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n487_), .B(KEYINPUT81), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n478_), .B1(new_n498_), .B2(new_n485_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n499_), .A2(new_n495_), .A3(new_n473_), .A4(new_n467_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n500_), .A3(KEYINPUT92), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n474_), .B(new_n502_), .C1(new_n490_), .C2(new_n496_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT4), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT93), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n497_), .A2(KEYINPUT4), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n506_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G57gat), .B(G85gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT95), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(new_n332_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n514_));
  INV_X1    g313(.A(G29gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n513_), .B(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n509_), .A2(new_n510_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n458_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n509_), .A2(new_n510_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n517_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n509_), .A2(new_n510_), .A3(new_n517_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(KEYINPUT99), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G71gat), .B(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G43gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT31), .ZN(new_n529_));
  INV_X1    g328(.A(new_n474_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(G15gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT30), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n534_), .A2(new_n399_), .A3(new_n411_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n411_), .B2(new_n399_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n412_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n534_), .A2(new_n399_), .A3(new_n411_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n474_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n529_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n529_), .A3(new_n541_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(KEYINPUT80), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT86), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n499_), .A2(new_n495_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT28), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n499_), .A2(new_n495_), .A3(new_n550_), .A4(new_n547_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G22gat), .B(G50gat), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n549_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n546_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n551_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT86), .A3(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n384_), .A2(new_n383_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n561_), .A2(new_n382_), .B1(new_n371_), .B2(new_n379_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n547_), .B1(new_n499_), .B2(new_n495_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G78gat), .B(G106gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT85), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT29), .B1(new_n490_), .B2(new_n496_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n386_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G228gat), .ZN(new_n570_));
  INV_X1    g369(.A(G233gat), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n566_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n565_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n386_), .A2(new_n568_), .A3(new_n567_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n555_), .B(new_n560_), .C1(new_n573_), .C2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT80), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n537_), .A2(new_n529_), .A3(new_n541_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n542_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT86), .B1(new_n558_), .B2(new_n559_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n572_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n575_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  AND4_X1   g384(.A1(new_n545_), .A2(new_n578_), .A3(new_n581_), .A4(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n543_), .A2(new_n544_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n578_), .B2(new_n585_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n520_), .B(new_n525_), .C1(new_n586_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n450_), .A2(new_n452_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n524_), .A2(KEYINPUT96), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n517_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n524_), .A2(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT96), .B1(new_n524_), .B2(new_n592_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n591_), .A2(new_n593_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n451_), .B2(KEYINPUT98), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n444_), .A2(new_n446_), .A3(new_n600_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n451_), .B2(new_n603_), .ZN(new_n604_));
  OAI22_X1  g403(.A1(new_n601_), .A2(new_n604_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n578_), .A2(new_n585_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n545_), .A2(new_n581_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n457_), .A2(new_n590_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n343_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G229gat), .A2(G233gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n343_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n298_), .A3(new_n294_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n343_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n616_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n614_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n622_), .B(new_n623_), .Z(new_n624_));
  AND3_X1   g423(.A1(new_n617_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n617_), .B2(new_n621_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n612_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n617_), .A2(new_n621_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n617_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(KEYINPUT76), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n611_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n357_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n520_), .A2(new_n525_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n332_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT38), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n324_), .A2(new_n327_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n611_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n355_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n625_), .A2(new_n626_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n279_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n635_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n640_), .B1(new_n648_), .B2(G1gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n639_), .B1(new_n649_), .B2(new_n636_), .ZN(G1324gat));
  INV_X1    g449(.A(new_n457_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n634_), .A2(new_n333_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n651_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  INV_X1    g458(.A(new_n647_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n609_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G15gat), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT102), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT102), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(KEYINPUT41), .A3(new_n664_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n634_), .A2(new_n532_), .A3(new_n609_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(G1326gat));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n647_), .B2(new_n608_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT42), .Z(new_n673_));
  NAND3_X1  g472(.A1(new_n634_), .A2(new_n671_), .A3(new_n608_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1327gat));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n611_), .B2(new_n331_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n328_), .A2(new_n330_), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n448_), .B(new_n589_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n610_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT43), .B(new_n678_), .C1(new_n679_), .C2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n279_), .A2(new_n645_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n677_), .A2(new_n644_), .A3(new_n682_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n678_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n355_), .B1(new_n687_), .B2(new_n676_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(KEYINPUT44), .A3(new_n683_), .A4(new_n682_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n686_), .A2(new_n689_), .A3(G29gat), .A4(new_n635_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n642_), .A2(new_n644_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n279_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n633_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n635_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n515_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n690_), .A2(new_n695_), .ZN(G1328gat));
  NOR3_X1   g495(.A1(new_n693_), .A2(G36gat), .A3(new_n457_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n686_), .A2(new_n689_), .A3(new_n651_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(KEYINPUT103), .A3(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n700_), .B2(G36gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n699_), .B(KEYINPUT46), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  INV_X1    g506(.A(new_n587_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n686_), .A2(new_n689_), .A3(G43gat), .A4(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n527_), .B1(new_n693_), .B2(new_n661_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g511(.A1(new_n686_), .A2(new_n689_), .A3(G50gat), .A4(new_n608_), .ZN(new_n713_));
  INV_X1    g512(.A(G50gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n693_), .B2(new_n607_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1331gat));
  NAND2_X1  g515(.A1(new_n630_), .A2(new_n631_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n611_), .A2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n277_), .A2(new_n278_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n356_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n635_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n719_), .B(KEYINPUT68), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n627_), .A2(new_n632_), .A3(new_n355_), .ZN(new_n725_));
  NOR4_X1   g524(.A1(new_n724_), .A2(new_n611_), .A3(new_n642_), .A4(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n635_), .B2(KEYINPUT104), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(KEYINPUT104), .B2(new_n727_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n723_), .B1(new_n726_), .B2(new_n729_), .ZN(G1332gat));
  INV_X1    g529(.A(G64gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n726_), .B2(new_n651_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT48), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n722_), .A2(new_n731_), .A3(new_n651_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n726_), .B2(new_n609_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT49), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n722_), .A2(new_n736_), .A3(new_n609_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  OR3_X1    g539(.A1(new_n721_), .A2(G78gat), .A3(new_n607_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n726_), .A2(new_n608_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G78gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT105), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n741_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1335gat));
  NOR4_X1   g549(.A1(new_n724_), .A2(new_n611_), .A3(new_n717_), .A4(new_n691_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n635_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n719_), .A2(new_n717_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n677_), .A2(new_n644_), .A3(new_n682_), .A4(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT106), .Z(new_n755_));
  NOR2_X1   g554(.A1(new_n694_), .A2(new_n209_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1336gat));
  AOI21_X1  g556(.A(G92gat), .B1(new_n751_), .B2(new_n651_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n457_), .A2(new_n210_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT107), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n755_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n751_), .A2(new_n708_), .A3(new_n204_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G99gat), .B1(new_n754_), .B2(new_n661_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g566(.A(G106gat), .B1(new_n754_), .B2(new_n607_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n751_), .A2(new_n205_), .A3(new_n608_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n770_), .B(new_n771_), .C1(new_n768_), .C2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT53), .ZN(G1339gat));
  XOR2_X1   g573(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n775_));
  NAND2_X1  g574(.A1(new_n613_), .A2(new_n616_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n613_), .A2(KEYINPUT114), .A3(new_n616_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n620_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n624_), .B1(new_n619_), .B2(new_n614_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n625_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n275_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n261_), .A2(KEYINPUT112), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n247_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n265_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n263_), .A2(new_n259_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n256_), .A2(KEYINPUT67), .A3(new_n202_), .A4(new_n257_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT55), .A3(new_n248_), .A4(new_n247_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n786_), .A2(new_n788_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n261_), .B2(new_n785_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n270_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n271_), .A2(new_n796_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT113), .B(new_n798_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n645_), .B2(new_n273_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n717_), .A2(KEYINPUT111), .A3(new_n272_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n784_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n775_), .B1(new_n808_), .B2(new_n642_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n805_), .A2(new_n806_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n800_), .A2(new_n799_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n802_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT57), .B(new_n641_), .C1(new_n812_), .C2(new_n784_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n793_), .A2(new_n794_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n815_), .A2(new_n798_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n782_), .A2(new_n272_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n814_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT58), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n820_), .A3(new_n678_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n809_), .A2(new_n813_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n644_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n725_), .A2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n627_), .A2(new_n632_), .A3(KEYINPUT110), .A4(new_n355_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n277_), .A3(new_n278_), .A4(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n827_), .B2(new_n678_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n277_), .A2(new_n278_), .A3(new_n826_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n331_), .A4(new_n825_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n823_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n457_), .A2(new_n635_), .A3(new_n588_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT116), .Z(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n822_), .B2(new_n644_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n837_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n717_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n837_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n813_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n809_), .A2(new_n821_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(KEYINPUT118), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n641_), .B1(new_n812_), .B2(new_n784_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n331_), .B1(KEYINPUT58), .B2(new_n819_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n850_), .A2(new_n775_), .B1(new_n818_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n355_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n846_), .B1(new_n855_), .B2(new_n832_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n839_), .B2(new_n840_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n627_), .B2(new_n632_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT119), .Z(new_n861_));
  AOI21_X1  g660(.A(new_n843_), .B1(new_n858_), .B2(new_n861_), .ZN(G1340gat));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n813_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n848_), .A2(KEYINPUT118), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n644_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n845_), .B1(new_n866_), .B2(new_n833_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n857_), .A2(new_n280_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n863_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n856_), .A2(KEYINPUT120), .A3(new_n280_), .A4(new_n857_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(G120gat), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n719_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n842_), .B(new_n873_), .C1(KEYINPUT60), .C2(new_n872_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1341gat));
  NAND3_X1  g674(.A1(new_n838_), .A2(new_n841_), .A3(new_n355_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n463_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT121), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(new_n879_), .A3(new_n463_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT122), .B(G127gat), .Z(new_n881_));
  NOR2_X1   g680(.A1(new_n644_), .A2(new_n881_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n878_), .A2(new_n880_), .B1(new_n858_), .B2(new_n882_), .ZN(G1342gat));
  AOI21_X1  g682(.A(G134gat), .B1(new_n842_), .B2(new_n642_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n678_), .A2(G134gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT123), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n858_), .B2(new_n886_), .ZN(G1343gat));
  INV_X1    g686(.A(new_n586_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n839_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n651_), .A2(new_n694_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n645_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n724_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(G148gat), .Z(G1345gat));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n355_), .A3(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n889_), .A2(new_n898_), .A3(new_n355_), .A4(new_n890_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  AND3_X1   g702(.A1(new_n889_), .A2(new_n678_), .A3(new_n890_), .ZN(new_n904_));
  INV_X1    g703(.A(G162gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n642_), .A2(new_n905_), .ZN(new_n906_));
  OAI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n891_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT125), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  OAI221_X1 g708(.A(new_n909_), .B1(new_n891_), .B2(new_n906_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1347gat));
  NOR3_X1   g710(.A1(new_n457_), .A2(new_n635_), .A3(new_n661_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n912_), .A2(new_n607_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n717_), .B(new_n913_), .C1(new_n855_), .C2(new_n832_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G169gat), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n387_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n917_), .B(new_n918_), .C1(new_n919_), .C2(new_n914_), .ZN(G1348gat));
  NAND2_X1  g719(.A1(new_n866_), .A2(new_n833_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n279_), .A3(new_n913_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n834_), .A2(KEYINPUT126), .A3(new_n607_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n839_), .B2(new_n608_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n923_), .A2(new_n912_), .A3(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n724_), .A2(new_n388_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n388_), .A2(new_n922_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  NAND2_X1  g727(.A1(new_n921_), .A2(new_n913_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n929_), .A2(new_n400_), .A3(new_n644_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G183gat), .B1(new_n926_), .B2(new_n355_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n929_), .B2(new_n331_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n642_), .A2(new_n404_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n929_), .B2(new_n934_), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n457_), .A2(new_n635_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n889_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n645_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n365_), .ZN(G1352gat));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n724_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n366_), .ZN(G1353gat));
  INV_X1    g740(.A(new_n937_), .ZN(new_n942_));
  AOI211_X1 g741(.A(KEYINPUT63), .B(G211gat), .C1(new_n942_), .C2(new_n355_), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT63), .B(G211gat), .Z(new_n944_));
  AND3_X1   g743(.A1(new_n942_), .A2(new_n355_), .A3(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n943_), .A2(new_n945_), .ZN(G1354gat));
  OR3_X1    g745(.A1(new_n937_), .A2(G218gat), .A3(new_n641_), .ZN(new_n947_));
  OAI21_X1  g746(.A(G218gat), .B1(new_n937_), .B2(new_n331_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1355gat));
endmodule


