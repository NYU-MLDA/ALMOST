//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n208_), .B2(KEYINPUT1), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(KEYINPUT86), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(KEYINPUT86), .B2(new_n209_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G141gat), .B(G148gat), .Z(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  INV_X1    g022(.A(new_n206_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n208_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n208_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT87), .A3(new_n206_), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n222_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n205_), .B1(new_n213_), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT4), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n205_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(KEYINPUT4), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G57gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n237_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n236_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(G183gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT25), .B1(new_n258_), .B2(KEYINPUT79), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(KEYINPUT25), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n257_), .B(new_n259_), .C1(new_n260_), .C2(KEYINPUT79), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G169gat), .A2(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT24), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n256_), .B(new_n261_), .C1(new_n255_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT80), .ZN(new_n265_));
  INV_X1    g064(.A(G169gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(KEYINPUT22), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n269_));
  INV_X1    g068(.A(G176gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(KEYINPUT22), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n272_), .A2(KEYINPUT81), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n252_), .B1(G183gat), .B2(G190gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT82), .B1(new_n274_), .B2(new_n250_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(KEYINPUT81), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n251_), .B(new_n252_), .C1(G183gat), .C2(G190gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n262_), .B1(new_n278_), .B2(KEYINPUT82), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n264_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n264_), .B(KEYINPUT83), .C1(new_n277_), .C2(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G43gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n284_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT84), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT30), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n288_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n205_), .B(KEYINPUT31), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n292_), .A2(KEYINPUT85), .A3(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n293_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n292_), .B2(KEYINPUT85), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n294_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G197gat), .B(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n302_), .A2(new_n303_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n301_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n301_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G197gat), .B(G204gat), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT21), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n314_), .B2(new_n304_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT90), .B1(new_n315_), .B2(new_n308_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n284_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT95), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  AOI21_X1  g122(.A(new_n255_), .B1(new_n263_), .B2(KEYINPUT96), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(KEYINPUT96), .B2(new_n263_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n257_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n256_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n262_), .B(KEYINPUT97), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n268_), .A2(G169gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n271_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n329_), .B(new_n278_), .C1(G176gat), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n315_), .A2(new_n308_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT20), .B(new_n323_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n319_), .A2(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n282_), .A2(new_n283_), .A3(new_n317_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n337_), .B(new_n342_), .C1(new_n346_), .C2(new_n323_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n342_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n323_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n335_), .B1(new_n284_), .B2(new_n318_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(KEYINPUT99), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n337_), .B1(new_n346_), .B2(new_n323_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT99), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n348_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n249_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n343_), .A2(new_n345_), .A3(new_n323_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n334_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT100), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n319_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n323_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n359_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT27), .B(new_n347_), .C1(new_n365_), .C2(new_n342_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n358_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT91), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n231_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n373_), .B1(new_n231_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n372_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n231_), .A2(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT28), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n375_), .A3(new_n371_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT29), .B1(new_n213_), .B2(new_n228_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n231_), .A2(new_n374_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT88), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT89), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n318_), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n383_), .A2(new_n334_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT93), .B1(new_n382_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT92), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n311_), .A2(new_n316_), .A3(new_n389_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(KEYINPUT88), .B2(new_n386_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n398_), .A2(new_n385_), .B1(new_n392_), .B2(new_n391_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n378_), .A2(new_n381_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT93), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n395_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n395_), .B2(new_n403_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n370_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n401_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n403_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n395_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n369_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n300_), .A2(new_n367_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n363_), .A2(new_n364_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n359_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n354_), .A2(new_n419_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n420_), .A2(new_n249_), .A3(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(KEYINPUT33), .B(new_n246_), .C1(new_n247_), .C2(new_n243_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n242_), .B1(new_n238_), .B2(new_n244_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n230_), .A2(new_n236_), .A3(new_n234_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n229_), .A2(new_n237_), .A3(new_n233_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(new_n242_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n425_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n423_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n356_), .B2(new_n352_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n412_), .B(new_n406_), .C1(new_n422_), .C2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n413_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n432_), .B(KEYINPUT101), .C1(new_n433_), .C2(new_n367_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n367_), .B1(new_n412_), .B2(new_n406_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT101), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n299_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT102), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n415_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT76), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT6), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT8), .ZN(new_n451_));
  INV_X1    g250(.A(G85gat), .ZN(new_n452_));
  INV_X1    g251(.A(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G85gat), .A2(G92gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n448_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT6), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(KEYINPUT66), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(KEYINPUT66), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n448_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n447_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT67), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n456_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n467_), .B2(new_n456_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n457_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT10), .B(G99gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT64), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n454_), .A2(new_n477_), .A3(KEYINPUT9), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n477_), .B1(new_n454_), .B2(KEYINPUT9), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n455_), .B1(new_n454_), .B2(KEYINPUT9), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n449_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT68), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n472_), .A2(new_n485_), .A3(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G29gat), .B(G36gat), .Z(new_n488_));
  XOR2_X1   g287(.A(G43gat), .B(G50gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G232gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT34), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(KEYINPUT35), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n482_), .B(KEYINPUT71), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n472_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n490_), .B(KEYINPUT15), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(KEYINPUT35), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n491_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n443_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G190gat), .B(G218gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n506_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  OAI221_X1 g310(.A(new_n443_), .B1(new_n511_), .B2(new_n507_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n514_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n515_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G71gat), .B(G78gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n521_), .B1(KEYINPUT11), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT69), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n532_), .B(new_n533_), .Z(new_n534_));
  XNOR2_X1  g333(.A(new_n526_), .B(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n535_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n535_), .A2(new_n541_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n520_), .A2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n472_), .A2(new_n485_), .A3(new_n482_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n485_), .B1(new_n472_), .B2(new_n482_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n526_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT70), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n487_), .A2(new_n552_), .A3(new_n526_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n526_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n484_), .A2(new_n554_), .A3(new_n486_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n551_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G230gat), .ZN(new_n557_));
  INV_X1    g356(.A(G233gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n526_), .A2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n555_), .A2(new_n562_), .B1(new_n496_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n559_), .B1(new_n487_), .B2(new_n526_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n560_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G120gat), .B(G148gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n560_), .A2(new_n567_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT75), .ZN(new_n586_));
  INV_X1    g385(.A(new_n490_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n532_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n532_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n532_), .B2(new_n497_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  MUX2_X1   g391(.A(new_n588_), .B(new_n591_), .S(new_n592_), .Z(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G169gat), .B(G197gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT78), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n593_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n586_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n442_), .A2(new_n547_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT103), .ZN(new_n603_));
  INV_X1    g402(.A(new_n430_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n352_), .A2(new_n356_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n418_), .A2(new_n419_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n604_), .A2(new_n605_), .B1(new_n606_), .B2(new_n421_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT101), .B1(new_n413_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n435_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n357_), .A2(new_n366_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n413_), .A2(new_n436_), .A3(new_n611_), .A4(new_n358_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n300_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT102), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n414_), .B1(new_n614_), .B2(new_n439_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n581_), .A2(new_n584_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n599_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n598_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n600_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n547_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n603_), .A2(KEYINPUT104), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT104), .B1(new_n603_), .B2(new_n623_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n202_), .B(new_n249_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n601_), .A2(new_n545_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n513_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n442_), .A2(KEYINPUT105), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n615_), .B2(new_n513_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n630_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n358_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n628_), .A2(new_n629_), .A3(new_n637_), .ZN(G1324gat));
  NOR2_X1   g437(.A1(new_n611_), .A2(G8gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n610_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(G8gat), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT39), .B(new_n528_), .C1(new_n635_), .C2(new_n610_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n640_), .B(KEYINPUT40), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  NAND2_X1  g448(.A1(new_n603_), .A2(new_n623_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n650_), .A2(G15gat), .A3(new_n300_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n635_), .A2(new_n299_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n652_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT41), .B1(new_n652_), .B2(G15gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n651_), .B1(new_n653_), .B2(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n635_), .A2(new_n413_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(G22gat), .ZN(new_n658_));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT42), .B(new_n659_), .C1(new_n635_), .C2(new_n413_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n413_), .A2(new_n659_), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n658_), .A2(new_n660_), .B1(new_n650_), .B2(new_n661_), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n631_), .A2(new_n545_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n621_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G29gat), .B1(new_n664_), .B2(new_n249_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n442_), .A2(new_n666_), .A3(new_n520_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n615_), .B2(new_n519_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n601_), .A2(new_n546_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n673_), .B(new_n670_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n249_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n665_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n675_), .B2(new_n610_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n664_), .A2(new_n679_), .A3(new_n610_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n680_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n681_), .B(KEYINPUT45), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n672_), .A2(new_n674_), .A3(new_n611_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n685_), .B(KEYINPUT46), .C1(new_n679_), .C2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1329gat));
  NAND2_X1  g487(.A1(new_n299_), .A2(G43gat), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n672_), .A2(new_n674_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G43gat), .B1(new_n664_), .B2(new_n299_), .ZN(new_n691_));
  OR3_X1    g490(.A1(new_n690_), .A2(KEYINPUT47), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT47), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n664_), .B2(new_n413_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n413_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n675_), .B2(new_n696_), .ZN(G1331gat));
  NOR2_X1   g496(.A1(new_n586_), .A2(new_n600_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n545_), .A3(new_n598_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(G57gat), .A3(new_n249_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(new_n703_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n615_), .A2(new_n618_), .A3(new_n698_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n547_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n249_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n704_), .A2(new_n705_), .A3(new_n709_), .ZN(G1332gat));
  INV_X1    g509(.A(G64gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n708_), .A2(new_n711_), .A3(new_n610_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n701_), .A2(new_n610_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G64gat), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT48), .B(new_n711_), .C1(new_n701_), .C2(new_n610_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1333gat));
  OR3_X1    g516(.A1(new_n707_), .A2(G71gat), .A3(new_n300_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n701_), .A2(new_n299_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G71gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G71gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1334gat));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n708_), .A2(new_n724_), .A3(new_n413_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n701_), .A2(new_n413_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G78gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT50), .B(new_n724_), .C1(new_n701_), .C2(new_n413_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1335gat));
  NAND2_X1  g529(.A1(new_n706_), .A2(new_n663_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n452_), .B1(new_n731_), .B2(new_n358_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT107), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n452_), .C1(new_n731_), .C2(new_n358_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n699_), .A2(new_n546_), .A3(new_n598_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(G85gat), .A3(new_n249_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n735_), .A3(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT108), .ZN(G1336gat));
  NAND2_X1  g539(.A1(new_n610_), .A2(G92gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT109), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n706_), .A2(new_n610_), .A3(new_n663_), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n737_), .A2(new_n742_), .B1(new_n743_), .B2(new_n453_), .ZN(G1337gat));
  INV_X1    g543(.A(G99gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n737_), .B2(new_n299_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n474_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n731_), .A2(new_n747_), .A3(new_n300_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n737_), .A2(new_n413_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G106gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT52), .B(new_n475_), .C1(new_n737_), .C2(new_n413_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n413_), .A2(new_n475_), .ZN(new_n755_));
  OAI22_X1  g554(.A1(new_n753_), .A2(new_n754_), .B1(new_n731_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  OAI221_X1 g557(.A(new_n758_), .B1(new_n731_), .B2(new_n755_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n598_), .A2(new_n545_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT110), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n519_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n765_), .B2(new_n585_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n764_), .A2(new_n616_), .A3(KEYINPUT54), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n574_), .A2(new_n618_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n496_), .A2(new_n564_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n548_), .A2(new_n549_), .A3(new_n526_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n561_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n550_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT112), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n567_), .A2(new_n779_), .A3(new_n772_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n565_), .A2(new_n566_), .A3(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n551_), .A2(new_n553_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n559_), .B1(new_n782_), .B2(new_n775_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .A4(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n576_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n770_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n591_), .A2(G229gat), .A3(G233gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n596_), .B1(new_n588_), .B2(new_n592_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT113), .Z(new_n793_));
  INV_X1    g592(.A(new_n596_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n593_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n578_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n631_), .B1(new_n789_), .B2(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n574_), .A2(new_n796_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n576_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n576_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n519_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT58), .B(new_n800_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n769_), .A2(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n770_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n797_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n631_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n807_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n768_), .B1(new_n812_), .B2(new_n546_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n611_), .A2(new_n249_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n300_), .A2(new_n814_), .A3(new_n413_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817_), .B2(new_n618_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n811_), .B1(new_n807_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n799_), .A2(new_n769_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n805_), .A2(new_n806_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n546_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n768_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT59), .B1(new_n813_), .B2(new_n816_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n618_), .A2(G113gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT115), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n818_), .B1(new_n831_), .B2(new_n833_), .ZN(G1340gat));
  NAND2_X1  g633(.A1(new_n803_), .A2(new_n804_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n835_), .A2(new_n520_), .A3(new_n806_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT57), .B1(new_n810_), .B2(new_n631_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT114), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n811_), .A3(new_n823_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n768_), .B1(new_n839_), .B2(new_n546_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n828_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n830_), .B(new_n699_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT117), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n829_), .A2(new_n844_), .A3(new_n699_), .A4(new_n830_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n845_), .A3(G120gat), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n698_), .A2(KEYINPUT60), .ZN(new_n847_));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  MUX2_X1   g647(.A(KEYINPUT60), .B(new_n847_), .S(new_n848_), .Z(new_n849_));
  NAND2_X1  g648(.A1(new_n817_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n846_), .A2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n817_), .A2(new_n854_), .A3(new_n545_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n829_), .A2(new_n545_), .A3(new_n830_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(new_n854_), .ZN(G1342gat));
  NAND4_X1  g657(.A1(new_n829_), .A2(G134gat), .A3(new_n520_), .A4(new_n830_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n813_), .A2(new_n631_), .A3(new_n816_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n860_), .A2(new_n861_), .A3(G134gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(G134gat), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n859_), .A2(new_n862_), .A3(new_n863_), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n300_), .A2(new_n413_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n814_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT119), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n813_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n618_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n699_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g671(.A(new_n868_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT120), .B1(new_n873_), .B2(new_n546_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n868_), .A2(new_n875_), .A3(new_n545_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n874_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1346gat));
  OR3_X1    g681(.A1(new_n873_), .A2(G162gat), .A3(new_n631_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G162gat), .B1(new_n873_), .B2(new_n519_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1347gat));
  NAND3_X1  g684(.A1(new_n299_), .A2(new_n358_), .A3(new_n610_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT121), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n413_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n827_), .A2(KEYINPUT125), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  INV_X1    g689(.A(new_n888_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n840_), .B2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n598_), .A2(new_n331_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n889_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n895_));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  OR3_X1    g695(.A1(new_n887_), .A2(new_n896_), .A3(new_n598_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n887_), .B2(new_n598_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n413_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n266_), .B1(new_n901_), .B2(KEYINPUT123), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n840_), .B2(new_n900_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n895_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n811_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n821_), .A2(new_n822_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(KEYINPUT114), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n545_), .B1(new_n908_), .B2(new_n823_), .ZN(new_n909_));
  OAI211_X1 g708(.A(KEYINPUT123), .B(new_n899_), .C1(new_n909_), .C2(new_n768_), .ZN(new_n910_));
  AND4_X1   g709(.A1(G169gat), .A2(new_n904_), .A3(new_n895_), .A4(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n894_), .B1(new_n905_), .B2(new_n911_), .ZN(G1348gat));
  INV_X1    g711(.A(new_n813_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n888_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n914_), .A2(new_n270_), .A3(new_n698_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n889_), .A2(new_n699_), .A3(new_n892_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n270_), .ZN(G1349gat));
  NOR2_X1   g716(.A1(new_n546_), .A2(new_n326_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n889_), .A2(new_n892_), .A3(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n258_), .B1(new_n914_), .B2(new_n546_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1350gat));
  NAND4_X1  g720(.A1(new_n889_), .A2(new_n892_), .A3(new_n513_), .A4(new_n257_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n889_), .A2(new_n520_), .A3(new_n892_), .ZN(new_n923_));
  INV_X1    g722(.A(G190gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n610_), .A2(new_n358_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n865_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n813_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n618_), .ZN(new_n930_));
  INV_X1    g729(.A(G197gat), .ZN(new_n931_));
  OR3_X1    g730(.A1(new_n930_), .A2(KEYINPUT126), .A3(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT126), .B1(new_n930_), .B2(new_n931_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n930_), .A2(new_n931_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n932_), .A2(new_n933_), .A3(new_n934_), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n929_), .A2(new_n699_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g736(.A1(new_n929_), .A2(new_n545_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT63), .B(G211gat), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941_));
  INV_X1    g740(.A(G211gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n938_), .A2(new_n941_), .A3(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n938_), .A2(KEYINPUT127), .A3(new_n941_), .A4(new_n942_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n940_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  INV_X1    g746(.A(new_n929_), .ZN(new_n948_));
  OR3_X1    g747(.A1(new_n948_), .A2(G218gat), .A3(new_n631_), .ZN(new_n949_));
  OAI21_X1  g748(.A(G218gat), .B1(new_n948_), .B2(new_n519_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1355gat));
endmodule


