//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n210_));
  INV_X1    g009(.A(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n207_), .B(new_n212_), .C1(new_n206_), .C2(new_n214_), .ZN(new_n215_));
  MUX2_X1   g014(.A(KEYINPUT23), .B(new_n210_), .S(new_n211_), .Z(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT85), .B(G176gat), .Z(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n213_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G71gat), .B(G99gat), .Z(new_n223_));
  XNOR2_X1  g022(.A(G15gat), .B(G43gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n222_), .B(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G127gat), .B(G134gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(G113gat), .B(G120gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n226_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT86), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT30), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT31), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n212_), .B1(G183gat), .B2(G190gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n219_), .B(KEYINPUT95), .ZN(new_n239_));
  INV_X1    g038(.A(new_n218_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n238_), .B(new_n213_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n206_), .A2(new_n205_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n216_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT94), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n213_), .A2(KEYINPUT93), .A3(KEYINPUT24), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n206_), .B1(new_n214_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n204_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n243_), .A2(KEYINPUT94), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n241_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n252_), .A2(G197gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(G197gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT21), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT92), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n253_), .B1(new_n257_), .B2(new_n254_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n257_), .B2(new_n254_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n255_), .B(new_n256_), .C1(new_n259_), .C2(KEYINPUT21), .ZN(new_n260_));
  INV_X1    g059(.A(new_n256_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(KEYINPUT21), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n251_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n222_), .A2(new_n263_), .ZN(new_n267_));
  OR3_X1    g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n251_), .A2(new_n263_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n269_), .B(KEYINPUT20), .C1(new_n263_), .C2(new_n222_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n272_), .A2(KEYINPUT97), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT97), .B1(new_n272_), .B2(new_n277_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n278_), .A2(KEYINPUT27), .A3(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n270_), .A2(new_n266_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n267_), .B1(new_n264_), .B2(KEYINPUT96), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n282_), .B1(KEYINPUT96), .B2(new_n264_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n283_), .B2(new_n266_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(new_n276_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n272_), .B(new_n276_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT27), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT89), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(KEYINPUT3), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n292_), .B(new_n297_), .C1(KEYINPUT3), .C2(new_n296_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n298_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n296_), .A2(KEYINPUT87), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(KEYINPUT87), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n299_), .B1(new_n300_), .B2(KEYINPUT1), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n299_), .A2(KEYINPUT1), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n310_));
  AOI211_X1 g109(.A(new_n303_), .B(new_n305_), .C1(new_n308_), .C2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n302_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(new_n229_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT4), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(new_n229_), .C1(new_n302_), .C2(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320_));
  INV_X1    g119(.A(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G57gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n313_), .A2(new_n318_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n319_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n319_), .B2(new_n325_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n302_), .A2(new_n311_), .A3(KEYINPUT29), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT28), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT90), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G228gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(G78gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G106gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n332_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n263_), .B1(new_n312_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT91), .Z(new_n341_));
  XOR2_X1   g140(.A(G22gat), .B(G50gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n338_), .A2(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n329_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n290_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n237_), .B1(new_n347_), .B2(KEYINPUT98), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n268_), .A2(new_n271_), .A3(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n328_), .B(new_n350_), .C1(new_n284_), .C2(new_n349_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n327_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n327_), .A2(new_n352_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n324_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n353_), .A2(new_n287_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n344_), .A2(new_n345_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT98), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n344_), .A2(new_n345_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n288_), .B1(new_n280_), .B2(new_n285_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n329_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n290_), .A2(new_n362_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n237_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n328_), .A2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n348_), .A2(new_n365_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT7), .ZN(new_n370_));
  INV_X1    g169(.A(G99gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n336_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G99gat), .A2(G106gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT65), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(KEYINPUT6), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(KEYINPUT65), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(KEYINPUT65), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(KEYINPUT6), .ZN(new_n382_));
  AND2_X1   g181(.A1(G99gat), .A2(G106gat), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n374_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G92gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n321_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G85gat), .A2(G92gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT67), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT8), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n372_), .A2(new_n373_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT8), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n390_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n394_), .A2(new_n395_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n387_), .A2(KEYINPUT9), .A3(new_n388_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n388_), .A2(KEYINPUT9), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT10), .B(G99gat), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n401_), .B(new_n402_), .C1(G106gat), .C2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT66), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n380_), .A2(new_n384_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n401_), .A2(new_n402_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n336_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n405_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n399_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT69), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n399_), .A2(new_n412_), .A3(KEYINPUT69), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT12), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G71gat), .B(G78gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(G57gat), .B(G64gat), .Z(new_n419_));
  INV_X1    g218(.A(KEYINPUT11), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT68), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G57gat), .B(G64gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(KEYINPUT11), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT68), .B1(new_n425_), .B2(new_n418_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n419_), .A2(new_n420_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n423_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n417_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n415_), .A2(new_n416_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n413_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n430_), .A2(new_n431_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n417_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n415_), .A2(KEYINPUT70), .A3(new_n416_), .A4(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G230gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT64), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n435_), .A2(new_n438_), .A3(new_n439_), .A4(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n437_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n436_), .A2(new_n437_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n441_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G120gat), .B(G148gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G176gat), .B(G204gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT72), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(new_n447_), .A3(new_n453_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT74), .Z(new_n461_));
  XNOR2_X1  g260(.A(G29gat), .B(G36gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT75), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT15), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467_));
  INV_X1    g266(.A(G1gat), .ZN(new_n468_));
  INV_X1    g267(.A(G8gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n473_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n465_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n465_), .B(new_n477_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n474_), .A2(new_n478_), .B1(new_n479_), .B2(new_n476_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G113gat), .B(G141gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT81), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n482_), .B(KEYINPUT82), .Z(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT83), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  OR3_X1    g285(.A1(new_n486_), .A2(new_n480_), .A3(new_n485_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n461_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n369_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n466_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n436_), .A2(new_n465_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G232gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT34), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n493_), .B(new_n494_), .C1(KEYINPUT35), .C2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(KEYINPUT35), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  XNOR2_X1  g298(.A(G190gat), .B(G218gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT76), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n499_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n503_), .B(KEYINPUT36), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n499_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n499_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n507_), .B(KEYINPUT77), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT37), .B1(new_n513_), .B2(new_n506_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n473_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n437_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT79), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(G183gat), .B(G211gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n519_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n518_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n524_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(KEYINPUT17), .B2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n518_), .A2(new_n526_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT80), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n515_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n492_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT99), .Z(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n468_), .A3(new_n328_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT38), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n531_), .ZN(new_n540_));
  NOR4_X1   g339(.A1(new_n369_), .A2(new_n491_), .A3(new_n508_), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(G1gat), .B1(new_n542_), .B2(new_n329_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n538_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n543_), .A3(new_n544_), .ZN(G1324gat));
  OAI21_X1  g344(.A(G8gat), .B1(new_n542_), .B2(new_n363_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT39), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n536_), .A2(new_n469_), .A3(new_n290_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(G1325gat));
  INV_X1    g350(.A(G15gat), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n541_), .B2(new_n237_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT101), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT41), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT41), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n536_), .A2(new_n552_), .A3(new_n237_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(G1326gat));
  INV_X1    g357(.A(G22gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n541_), .B2(new_n362_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT42), .Z(new_n561_));
  NAND3_X1  g360(.A1(new_n536_), .A2(new_n559_), .A3(new_n362_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(G1327gat));
  AND2_X1   g362(.A1(new_n508_), .A2(new_n533_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n492_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(G29gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n328_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT102), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n348_), .A2(new_n365_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n366_), .A2(new_n368_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n515_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT43), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n532_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(KEYINPUT43), .A3(new_n515_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(KEYINPUT44), .A3(new_n490_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n510_), .A2(new_n514_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n574_), .B1(new_n369_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n576_), .A2(new_n579_), .A3(new_n533_), .A4(new_n490_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT44), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n328_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n569_), .B1(new_n584_), .B2(G29gat), .ZN(new_n585_));
  AOI211_X1 g384(.A(KEYINPUT102), .B(new_n567_), .C1(new_n583_), .C2(new_n328_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n568_), .B1(new_n585_), .B2(new_n586_), .ZN(G1328gat));
  NOR3_X1   g386(.A1(new_n565_), .A2(G36gat), .A3(new_n363_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT45), .Z(new_n589_));
  NAND3_X1  g388(.A1(new_n577_), .A2(new_n582_), .A3(new_n290_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT103), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G36gat), .B1(new_n590_), .B2(new_n591_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI221_X1 g395(.A(new_n589_), .B1(KEYINPUT104), .B2(KEYINPUT46), .C1(new_n592_), .C2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(G1329gat));
  NOR3_X1   g397(.A1(new_n565_), .A2(G43gat), .A3(new_n367_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n583_), .A2(new_n237_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n600_), .B2(G43gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n601_), .B(new_n603_), .ZN(G1330gat));
  AOI21_X1  g403(.A(G50gat), .B1(new_n566_), .B2(new_n362_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n362_), .A2(G50gat), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n583_), .B2(new_n606_), .ZN(G1331gat));
  INV_X1    g406(.A(new_n489_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n461_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n369_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(new_n534_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G57gat), .B1(new_n611_), .B2(new_n328_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n532_), .A2(new_n489_), .ZN(new_n613_));
  NOR4_X1   g412(.A1(new_n369_), .A2(new_n508_), .A3(new_n609_), .A4(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(G57gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n328_), .B2(KEYINPUT106), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(KEYINPUT106), .B2(new_n615_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n612_), .B1(new_n614_), .B2(new_n617_), .ZN(G1332gat));
  INV_X1    g417(.A(new_n614_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G64gat), .B1(new_n619_), .B2(new_n363_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT48), .ZN(new_n621_));
  INV_X1    g420(.A(G64gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n611_), .A2(new_n622_), .A3(new_n290_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT107), .ZN(G1333gat));
  INV_X1    g424(.A(G71gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n614_), .B2(new_n237_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT49), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n611_), .A2(new_n626_), .A3(new_n237_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1334gat));
  AOI21_X1  g429(.A(new_n334_), .B1(new_n614_), .B2(new_n362_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT50), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n611_), .A2(new_n334_), .A3(new_n362_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1335gat));
  NOR2_X1   g433(.A1(new_n609_), .A2(new_n608_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n576_), .A2(new_n579_), .A3(new_n533_), .A4(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G85gat), .B1(new_n636_), .B2(new_n329_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n610_), .A2(new_n564_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1336gat));
  OAI21_X1  g439(.A(G92gat), .B1(new_n636_), .B2(new_n363_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n386_), .A3(new_n290_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1337gat));
  OAI21_X1  g442(.A(G99gat), .B1(new_n636_), .B2(new_n367_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n638_), .A2(new_n408_), .A3(new_n237_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT51), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(KEYINPUT108), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n646_), .B(new_n648_), .ZN(G1338gat));
  NAND3_X1  g448(.A1(new_n638_), .A2(new_n336_), .A3(new_n362_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G106gat), .B1(new_n636_), .B2(new_n359_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT109), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT52), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT109), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n654_), .B(G106gat), .C1(new_n636_), .C2(new_n359_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n652_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n653_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n650_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n650_), .B(new_n659_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1339gat));
  INV_X1    g462(.A(KEYINPUT111), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n613_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n532_), .A2(new_n489_), .A3(KEYINPUT111), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n578_), .A2(new_n665_), .A3(new_n460_), .A4(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT54), .Z(new_n668_));
  INV_X1    g467(.A(KEYINPUT57), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n508_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n475_), .B1(new_n465_), .B2(new_n477_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n474_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n485_), .B1(new_n479_), .B2(new_n475_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n672_), .A2(new_n673_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n457_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n608_), .A2(new_n456_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n435_), .A2(new_n444_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n441_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT55), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n443_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n439_), .A2(new_n438_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n681_), .A2(KEYINPUT55), .A3(new_n435_), .A4(new_n442_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(KEYINPUT56), .A3(new_n454_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT113), .B(KEYINPUT56), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n454_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT112), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n690_), .A3(new_n454_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n687_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT114), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n685_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n683_), .A2(new_n690_), .A3(new_n454_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n690_), .B1(new_n683_), .B2(new_n454_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n686_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT114), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n676_), .B1(new_n694_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT115), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n675_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n676_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n684_), .B1(new_n697_), .B2(KEYINPUT114), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n689_), .A2(new_n691_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n693_), .B1(new_n704_), .B2(new_n686_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n700_), .B(new_n702_), .C1(new_n703_), .C2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n670_), .B1(new_n701_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT58), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT56), .B1(new_n683_), .B2(new_n454_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n456_), .B(new_n674_), .C1(new_n685_), .C2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n711_), .B2(KEYINPUT117), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT116), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT117), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n515_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n712_), .A2(new_n714_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n675_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n702_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(KEYINPUT115), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n508_), .B1(new_n720_), .B2(new_n706_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n708_), .B(new_n717_), .C1(new_n721_), .C2(KEYINPUT57), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n668_), .B1(new_n722_), .B2(new_n540_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n366_), .A2(new_n328_), .A3(new_n237_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT59), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT59), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n701_), .A2(new_n707_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n669_), .B1(new_n727_), .B2(new_n508_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n715_), .A2(new_n716_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n720_), .A2(new_n706_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n670_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n532_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n726_), .B1(new_n732_), .B2(new_n668_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n725_), .A2(KEYINPUT119), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT119), .B1(new_n725_), .B2(new_n733_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n489_), .ZN(new_n736_));
  INV_X1    g535(.A(G113gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n724_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n531_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT118), .B(new_n740_), .C1(new_n741_), .C2(new_n668_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n608_), .A2(new_n737_), .ZN(new_n744_));
  OAI22_X1  g543(.A1(new_n736_), .A2(new_n737_), .B1(new_n743_), .B2(new_n744_), .ZN(G1340gat));
  NAND3_X1  g544(.A1(new_n725_), .A2(new_n461_), .A3(new_n733_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G120gat), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT60), .ZN(new_n748_));
  AOI21_X1  g547(.A(G120gat), .B1(new_n461_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n748_), .B2(G120gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n742_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n751_), .ZN(G1341gat));
  INV_X1    g551(.A(G127gat), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n540_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n734_), .A2(new_n735_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n739_), .A2(new_n742_), .A3(new_n532_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n753_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT120), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n735_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n725_), .A2(KEYINPUT119), .A3(new_n733_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n754_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT120), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n758_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n760_), .A2(new_n765_), .ZN(G1342gat));
  NOR3_X1   g565(.A1(new_n734_), .A2(new_n735_), .A3(new_n578_), .ZN(new_n767_));
  INV_X1    g566(.A(G134gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n508_), .A2(new_n768_), .ZN(new_n769_));
  OAI22_X1  g568(.A1(new_n767_), .A2(new_n768_), .B1(new_n743_), .B2(new_n769_), .ZN(G1343gat));
  INV_X1    g569(.A(new_n723_), .ZN(new_n771_));
  NOR4_X1   g570(.A1(new_n290_), .A2(new_n359_), .A3(new_n329_), .A4(new_n237_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n489_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(new_n294_), .ZN(G1344gat));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n609_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT121), .B(G148gat), .Z(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(G1345gat));
  INV_X1    g577(.A(new_n773_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT122), .A3(new_n532_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT122), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n773_), .B2(new_n533_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT61), .B(G155gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(G1346gat));
  INV_X1    g584(.A(G162gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n779_), .A2(new_n786_), .A3(new_n508_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G162gat), .B1(new_n773_), .B2(new_n578_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT123), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n787_), .A2(KEYINPUT123), .A3(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1347gat));
  NOR2_X1   g592(.A1(new_n732_), .A2(new_n668_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n290_), .A2(new_n368_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(new_n362_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n608_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G169gat), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n799_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(G169gat), .A3(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n800_), .B(new_n802_), .C1(new_n239_), .C2(new_n797_), .ZN(G1348gat));
  NAND2_X1  g602(.A1(new_n771_), .A2(new_n359_), .ZN(new_n804_));
  INV_X1    g603(.A(G176gat), .ZN(new_n805_));
  NOR4_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n609_), .A4(new_n795_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n240_), .B1(new_n796_), .B2(new_n461_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT125), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(KEYINPUT125), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n806_), .B1(new_n808_), .B2(new_n809_), .ZN(G1349gat));
  OR3_X1    g609(.A1(new_n804_), .A2(new_n533_), .A3(new_n795_), .ZN(new_n811_));
  INV_X1    g610(.A(G183gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n540_), .A2(new_n202_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n811_), .A2(new_n812_), .B1(new_n796_), .B2(new_n813_), .ZN(G1350gat));
  NAND2_X1  g613(.A1(new_n796_), .A2(new_n515_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(G190gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n796_), .A2(new_n508_), .A3(new_n203_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1351gat));
  NAND3_X1  g617(.A1(new_n362_), .A2(new_n329_), .A3(new_n367_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n723_), .A2(new_n363_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n608_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G197gat), .ZN(G1352gat));
  OAI211_X1 g621(.A(new_n820_), .B(new_n461_), .C1(KEYINPUT126), .C2(new_n252_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n252_), .A2(KEYINPUT126), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT127), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n823_), .B(new_n825_), .ZN(G1353gat));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n531_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n828_));
  AND2_X1   g627(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n827_), .B2(new_n828_), .ZN(G1354gat));
  INV_X1    g630(.A(G218gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n832_), .A3(new_n508_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n820_), .A2(new_n515_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1355gat));
endmodule


