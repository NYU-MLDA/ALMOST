//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(G228gat), .ZN(new_n202_));
  INV_X1    g001(.A(G233gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT92), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT92), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G78gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT94), .A2(G204gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT94), .A2(G204gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(G197gat), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(KEYINPUT95), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT95), .B1(new_n210_), .B2(new_n212_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT96), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT95), .ZN(new_n220_));
  INV_X1    g019(.A(G197gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n209_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT94), .A2(G204gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n224_), .B2(new_n211_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT96), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n219_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G211gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G218gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(G218gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n208_), .A2(new_n209_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n221_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n215_), .B1(G197gat), .B2(G204gat), .ZN(new_n234_));
  AOI211_X1 g033(.A(new_n230_), .B(new_n231_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n215_), .B1(new_n224_), .B2(new_n211_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n228_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  OR3_X1    g039(.A1(new_n240_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT89), .B1(new_n240_), .B2(KEYINPUT1), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT88), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT88), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(G155gat), .B2(G162gat), .ZN(new_n247_));
  AOI22_X1  g046(.A1(new_n245_), .A2(new_n247_), .B1(KEYINPUT1), .B2(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT87), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(KEYINPUT87), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n249_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n250_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT91), .B1(KEYINPUT90), .B2(KEYINPUT3), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(new_n255_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n252_), .A2(new_n260_), .A3(new_n253_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n255_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n245_), .A2(new_n247_), .B1(G155gat), .B2(G162gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n239_), .B1(new_n259_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT93), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n238_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n219_), .A2(new_n227_), .B1(new_n236_), .B2(new_n235_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT93), .B1(new_n275_), .B2(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n259_), .A2(new_n270_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT28), .B1(new_n277_), .B2(KEYINPUT29), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n258_), .A2(new_n249_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n239_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n274_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G22gat), .B(G50gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n282_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n273_), .B1(new_n238_), .B2(new_n272_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n275_), .A2(new_n271_), .A3(KEYINPUT93), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n274_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n207_), .B1(new_n287_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT97), .B(G106gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n286_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n285_), .A3(new_n292_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n207_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G8gat), .B(G36gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT18), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n306_));
  INV_X1    g105(.A(G169gat), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT23), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G169gat), .B(G176gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n309_), .B(new_n311_), .C1(new_n312_), .C2(new_n306_), .ZN(new_n313_));
  INV_X1    g112(.A(G183gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT25), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G183gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT98), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(G190gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n313_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n310_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n323_), .B(new_n324_), .C1(G183gat), .C2(G190gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n326_));
  OR3_X1    g125(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n321_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n275_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n311_), .B(new_n333_), .C1(new_n332_), .C2(new_n312_), .ZN(new_n334_));
  INV_X1    g133(.A(G190gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT83), .B1(new_n335_), .B2(KEYINPUT26), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(new_n335_), .A3(KEYINPUT26), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT83), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT26), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(G190gat), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n336_), .A2(new_n338_), .A3(new_n341_), .A4(new_n317_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n316_), .B2(G183gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n314_), .A2(KEYINPUT81), .A3(KEYINPUT25), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n340_), .A2(G190gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n344_), .B(new_n345_), .C1(new_n346_), .C2(new_n337_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n328_), .B1(new_n334_), .B2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n238_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n331_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n330_), .B2(new_n275_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n238_), .A2(new_n349_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT32), .B(new_n305_), .C1(new_n353_), .C2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n331_), .B2(new_n350_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G120gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n367_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT84), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n277_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n370_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n259_), .A2(new_n270_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n365_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT100), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n374_), .B2(KEYINPUT4), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(KEYINPUT4), .A3(new_n376_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n277_), .A2(KEYINPUT100), .A3(new_n373_), .A4(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n383_), .B2(new_n365_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G1gat), .B(G29gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G57gat), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  AOI211_X1 g190(.A(new_n389_), .B(new_n377_), .C1(new_n383_), .C2(new_n365_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n359_), .B(new_n363_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n383_), .A2(new_n365_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT33), .B(new_n389_), .C1(new_n394_), .C2(new_n377_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n384_), .B2(new_n390_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n360_), .A2(new_n361_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n304_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n374_), .A2(new_n376_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n364_), .B1(new_n401_), .B2(KEYINPUT102), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(KEYINPUT102), .B2(new_n401_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n403_), .B(new_n390_), .C1(new_n365_), .C2(new_n383_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n360_), .A2(new_n305_), .A3(new_n361_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n400_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n393_), .B1(new_n398_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n295_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n298_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n349_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(G15gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT30), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n414_), .B(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(KEYINPUT85), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n373_), .B(KEYINPUT31), .Z(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n419_), .B(KEYINPUT85), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  AND4_X1   g223(.A1(new_n300_), .A2(new_n407_), .A3(new_n411_), .A4(new_n424_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n409_), .A2(new_n410_), .A3(new_n408_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n295_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n421_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n421_), .B2(new_n420_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n411_), .A3(new_n300_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n400_), .A2(new_n405_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT27), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n304_), .B1(new_n353_), .B2(new_n358_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT27), .A3(new_n405_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n391_), .A2(new_n392_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n425_), .B1(new_n432_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G113gat), .B(G141gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT79), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G169gat), .B(G197gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT74), .B(G15gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G22gat), .ZN(new_n448_));
  INV_X1    g247(.A(G1gat), .ZN(new_n449_));
  INV_X1    g248(.A(G8gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT14), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G1gat), .B(G8gat), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n452_), .B(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G29gat), .B(G36gat), .Z(new_n456_));
  XOR2_X1   g255(.A(G43gat), .B(G50gat), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n452_), .B(new_n453_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n458_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n462_), .A3(KEYINPUT77), .ZN(new_n463_));
  OR3_X1    g262(.A1(new_n461_), .A2(KEYINPUT77), .A3(new_n458_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G229gat), .A2(G233gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n458_), .B(KEYINPUT15), .Z(new_n468_));
  OR2_X1    g267(.A1(new_n468_), .A2(new_n461_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n465_), .A3(new_n462_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n446_), .B1(new_n471_), .B2(KEYINPUT78), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(KEYINPUT78), .B2(new_n471_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n470_), .A3(new_n446_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT80), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n467_), .A2(KEYINPUT80), .A3(new_n470_), .A4(new_n446_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n442_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT66), .ZN(new_n483_));
  AND3_X1   g282(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G85gat), .A2(G92gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT67), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n483_), .B(new_n486_), .C1(KEYINPUT67), .C2(new_n484_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT6), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n488_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(KEYINPUT6), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT68), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT10), .B(G99gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT65), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n487_), .B(new_n498_), .C1(G106gat), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G85gat), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(new_n485_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n506_));
  OR2_X1    g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT69), .ZN(new_n509_));
  NOR4_X1   g308(.A1(new_n509_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT7), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT69), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n508_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n497_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n494_), .A2(new_n495_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n517_), .B(new_n508_), .C1(new_n510_), .C2(new_n513_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n505_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n515_), .B1(new_n520_), .B2(KEYINPUT70), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n509_), .B1(new_n507_), .B2(KEYINPUT7), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(KEYINPUT69), .A3(new_n512_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n494_), .A2(new_n495_), .B1(new_n507_), .B2(KEYINPUT7), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n505_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n516_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n501_), .B1(new_n521_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n468_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n532_), .A2(KEYINPUT35), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n520_), .A2(KEYINPUT70), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n527_), .B1(new_n526_), .B2(new_n516_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n515_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n459_), .A3(new_n501_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT73), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n530_), .A2(new_n540_), .A3(new_n537_), .A4(new_n533_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n530_), .A2(new_n537_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n532_), .A2(KEYINPUT35), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n533_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n539_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G134gat), .B(G162gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n538_), .A2(KEYINPUT73), .B1(new_n542_), .B2(new_n544_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n554_), .A2(new_n550_), .A3(new_n549_), .A4(new_n541_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT64), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(KEYINPUT11), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n564_));
  INV_X1    g363(.A(new_n562_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n563_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n568_), .B(new_n501_), .C1(new_n521_), .C2(new_n528_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(new_n536_), .B2(new_n501_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n560_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(KEYINPUT71), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n574_), .B(new_n563_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(KEYINPUT12), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n529_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n571_), .B2(KEYINPUT12), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n569_), .A2(new_n559_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n572_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G120gat), .B(G148gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT13), .B1(new_n587_), .B2(new_n588_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT17), .ZN(new_n599_));
  INV_X1    g398(.A(new_n568_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n461_), .B(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n599_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n602_), .B2(new_n601_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(KEYINPUT71), .A3(KEYINPUT17), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT76), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n557_), .A2(new_n593_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n481_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n613_), .A2(G1gat), .A3(new_n439_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(KEYINPUT38), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT103), .Z(new_n616_));
  AND2_X1   g415(.A1(new_n553_), .A2(new_n555_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n442_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n593_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n480_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n618_), .A2(new_n610_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n439_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n449_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(KEYINPUT38), .B2(new_n614_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n616_), .A2(new_n624_), .ZN(G1324gat));
  NAND2_X1  g424(.A1(new_n435_), .A2(new_n437_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n450_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n626_), .A2(new_n450_), .ZN(new_n633_));
  OAI22_X1  g432(.A1(new_n631_), .A2(new_n632_), .B1(new_n613_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  AOI21_X1  g435(.A(new_n416_), .B1(new_n621_), .B2(new_n430_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n430_), .A2(new_n416_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n613_), .B2(new_n639_), .ZN(G1326gat));
  NOR2_X1   g439(.A1(new_n426_), .A2(new_n427_), .ZN(new_n641_));
  OR3_X1    g440(.A1(new_n613_), .A2(G22gat), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n621_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(G22gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n644_), .B2(G22gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n642_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT105), .ZN(G1327gat));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n442_), .B2(new_n557_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n556_), .B(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n440_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT43), .B(new_n654_), .C1(new_n655_), .C2(new_n425_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n652_), .A2(new_n609_), .A3(new_n620_), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n655_), .B2(new_n425_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n610_), .B1(new_n660_), .B2(new_n651_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n620_), .A4(new_n656_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n622_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G29gat), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n610_), .A2(new_n556_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n481_), .A2(new_n593_), .A3(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n439_), .A2(G29gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  OR2_X1    g467(.A1(new_n438_), .A2(G36gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT45), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n659_), .A2(new_n626_), .A3(new_n662_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT106), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n659_), .A2(new_n674_), .A3(new_n662_), .A4(new_n626_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G36gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n671_), .B(KEYINPUT46), .C1(new_n673_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  INV_X1    g480(.A(G43gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n666_), .B2(new_n424_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT107), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n659_), .A2(G43gat), .A3(new_n662_), .A4(new_n430_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g486(.A1(new_n659_), .A2(G50gat), .A3(new_n662_), .A4(new_n643_), .ZN(new_n688_));
  INV_X1    g487(.A(G50gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n666_), .B2(new_n641_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n442_), .A2(new_n479_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n654_), .A2(new_n609_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n619_), .ZN(new_n694_));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n622_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n593_), .A2(new_n479_), .A3(new_n609_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n618_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n439_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n694_), .A2(new_n701_), .A3(new_n626_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G64gat), .B1(new_n698_), .B2(new_n438_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n703_), .A2(new_n705_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n702_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g509(.A(G71gat), .B1(new_n698_), .B2(new_n424_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT49), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n424_), .A2(G71gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT110), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n694_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1334gat));
  OAI21_X1  g515(.A(G78gat), .B1(new_n698_), .B2(new_n641_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(G78gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n694_), .A2(new_n720_), .A3(new_n643_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1335gat));
  NOR2_X1   g521(.A1(new_n593_), .A2(new_n479_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n661_), .A2(new_n656_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n439_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n692_), .A2(new_n619_), .A3(new_n665_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n502_), .A3(new_n622_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1336gat));
  OAI21_X1  g527(.A(G92gat), .B1(new_n724_), .B2(new_n438_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n503_), .A3(new_n626_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1337gat));
  OAI21_X1  g530(.A(G99gat), .B1(new_n724_), .B2(new_n424_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n500_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n726_), .A2(new_n430_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g535(.A(G106gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n726_), .A2(new_n737_), .A3(new_n643_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n661_), .A2(new_n643_), .A3(new_n656_), .A4(new_n723_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(G106gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G106gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g543(.A(new_n431_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n626_), .A2(new_n439_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT12), .B1(new_n529_), .B2(new_n600_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n576_), .B1(new_n536_), .B2(new_n501_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n750_), .A2(new_n580_), .A3(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n578_), .B(new_n569_), .C1(new_n571_), .C2(KEYINPUT12), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n752_), .A2(KEYINPUT55), .B1(new_n560_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT112), .B1(new_n752_), .B2(KEYINPUT55), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n756_), .B(new_n757_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT56), .A3(new_n586_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT114), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n586_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(KEYINPUT114), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(new_n586_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n587_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n465_), .B1(new_n461_), .B2(new_n458_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n446_), .B1(new_n469_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n589_), .A2(new_n478_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n749_), .B1(new_n776_), .B2(new_n556_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n775_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n556_), .A2(KEYINPUT57), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n478_), .A2(new_n587_), .A3(new_n774_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n760_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n586_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n781_), .B(KEYINPUT58), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n654_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n762_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n760_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT58), .B1(new_n788_), .B2(new_n781_), .ZN(new_n789_));
  OAI22_X1  g588(.A1(new_n779_), .A2(new_n780_), .B1(new_n785_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n609_), .B1(new_n777_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT54), .B1(new_n611_), .B2(new_n479_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n693_), .A2(new_n793_), .A3(new_n480_), .A4(new_n593_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n747_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  INV_X1    g597(.A(new_n780_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n776_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n748_), .B1(new_n779_), .B2(new_n617_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n478_), .A2(new_n587_), .A3(new_n774_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n787_), .B2(new_n760_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n803_), .A2(KEYINPUT58), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n557_), .B1(new_n803_), .B2(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(new_n801_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n795_), .B1(new_n807_), .B2(new_n609_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n747_), .A2(KEYINPUT116), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n747_), .A2(KEYINPUT116), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n798_), .A3(new_n810_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n797_), .A2(new_n798_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n480_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n747_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(new_n776_), .A2(new_n799_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n610_), .B1(new_n815_), .B2(new_n801_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n814_), .B1(new_n816_), .B2(new_n795_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n480_), .A2(G113gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n813_), .B1(new_n817_), .B2(new_n818_), .ZN(G1340gat));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n811_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n817_), .B2(KEYINPUT59), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n823_), .B2(new_n619_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT117), .B1(new_n821_), .B2(KEYINPUT60), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n797_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n820_), .B1(new_n824_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G120gat), .B1(new_n812_), .B2(new_n593_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(KEYINPUT118), .A3(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1341gat));
  OAI21_X1  g634(.A(G127gat), .B1(new_n812_), .B2(new_n609_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n609_), .A2(G127gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n817_), .B2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n797_), .B2(new_n617_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n840_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT120), .B(G134gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n557_), .A2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n841_), .A2(new_n842_), .B1(new_n823_), .B2(new_n844_), .ZN(G1343gat));
  NAND2_X1  g644(.A1(new_n791_), .A2(new_n796_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n428_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n746_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n480_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n593_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT121), .B(G148gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1345gat));
  NOR2_X1   g652(.A1(new_n848_), .A2(new_n609_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n854_), .B(new_n855_), .Z(G1346gat));
  OAI21_X1  g655(.A(G162gat), .B1(new_n848_), .B2(new_n557_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n556_), .A2(G162gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n848_), .B2(new_n858_), .ZN(G1347gat));
  NOR2_X1   g658(.A1(new_n438_), .A2(new_n622_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n430_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n480_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT122), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n643_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n307_), .B1(new_n846_), .B2(new_n864_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT62), .Z(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n861_), .A2(new_n643_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n808_), .B2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n846_), .A2(KEYINPUT123), .A3(new_n868_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT22), .B(G169gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n479_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n866_), .A2(new_n874_), .ZN(G1348gat));
  NOR3_X1   g674(.A1(new_n808_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT123), .B1(new_n846_), .B2(new_n868_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n619_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n308_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n593_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT124), .B1(new_n881_), .B2(G176gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n808_), .A2(new_n869_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n593_), .A2(new_n308_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n880_), .A2(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  AOI21_X1  g684(.A(G183gat), .B1(new_n883_), .B2(new_n610_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n609_), .A2(new_n319_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n872_), .B2(new_n887_), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n872_), .A2(new_n320_), .A3(new_n617_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n557_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n335_), .B2(new_n890_), .ZN(G1351gat));
  NAND3_X1  g690(.A1(new_n846_), .A2(new_n847_), .A3(new_n860_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n480_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n221_), .ZN(G1352gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n593_), .ZN(new_n895_));
  MUX2_X1   g694(.A(G204gat), .B(new_n232_), .S(new_n895_), .Z(G1353gat));
  AND3_X1   g695(.A1(new_n846_), .A2(new_n847_), .A3(new_n860_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n609_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n900_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n898_), .B1(new_n892_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n901_), .A2(new_n905_), .A3(new_n903_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1354gat));
  AND3_X1   g708(.A1(new_n897_), .A2(G218gat), .A3(new_n654_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n892_), .A2(new_n556_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n911_), .A2(KEYINPUT127), .ZN(new_n912_));
  AOI21_X1  g711(.A(G218gat), .B1(new_n911_), .B2(KEYINPUT127), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n912_), .B2(new_n913_), .ZN(G1355gat));
endmodule


