//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203_));
  XOR2_X1   g002(.A(G113gat), .B(G120gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT31), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT91), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n206_), .B2(new_n205_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(G183gat), .B2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n211_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(KEYINPUT88), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(new_n212_), .A3(G183gat), .A4(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n213_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT24), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT87), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  INV_X1    g032(.A(G183gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT25), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT86), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G183gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT86), .B1(new_n235_), .B2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n230_), .B(new_n232_), .C1(new_n237_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n229_), .A2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n235_), .A2(new_n239_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n233_), .B(new_n236_), .C1(new_n243_), .C2(KEYINPUT86), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n230_), .B1(new_n244_), .B2(new_n232_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n220_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G15gat), .B(G43gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT90), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n246_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G227gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G71gat), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n252_), .A2(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n210_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n251_), .B(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n209_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT101), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT100), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G141gat), .ZN(new_n271_));
  INV_X1    g070(.A(G148gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT95), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT3), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n275_), .A2(new_n271_), .A3(new_n272_), .A4(KEYINPUT95), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n270_), .A2(new_n274_), .A3(new_n276_), .A4(new_n277_), .ZN(new_n278_));
  NOR3_X1   g077(.A1(KEYINPUT94), .A2(G155gat), .A3(G162gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT94), .B1(G155gat), .B2(G162gat), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n280_), .A2(new_n281_), .B1(G155gat), .B2(G162gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT93), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT93), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(G141gat), .B2(G148gat), .ZN(new_n285_));
  AND4_X1   g084(.A1(new_n267_), .A2(new_n283_), .A3(new_n285_), .A4(new_n269_), .ZN(new_n286_));
  INV_X1    g085(.A(G155gat), .ZN(new_n287_));
  INV_X1    g086(.A(G162gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT1), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(G155gat), .A3(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n281_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n289_), .B(new_n291_), .C1(new_n292_), .C2(new_n279_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n278_), .A2(new_n282_), .B1(new_n286_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n264_), .B1(new_n294_), .B2(new_n205_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n278_), .A2(new_n282_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n286_), .A2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n203_), .B(new_n204_), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n264_), .A3(new_n299_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n263_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(KEYINPUT4), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n262_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n262_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n306_), .A3(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G85gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT0), .B(G57gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n305_), .A2(new_n314_), .A3(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n294_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT28), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT97), .B1(new_n321_), .B2(G197gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT97), .ZN(new_n323_));
  INV_X1    g122(.A(G197gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(G204gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(G197gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT21), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT96), .B1(new_n321_), .B2(G197gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT96), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n324_), .A3(G204gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n333_), .A3(new_n326_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n330_), .B1(new_n334_), .B2(KEYINPUT21), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n329_), .A2(new_n336_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n328_), .A2(new_n335_), .B1(new_n327_), .B2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(KEYINPUT29), .B2(new_n298_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n320_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G78gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G106gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G22gat), .B(G50gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n340_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n328_), .A2(new_n335_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n337_), .A2(new_n327_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n228_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT26), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G190gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n235_), .A2(new_n239_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n362_), .A2(KEYINPUT98), .A3(new_n232_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT98), .B1(new_n362_), .B2(new_n232_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n357_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n219_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n217_), .A2(KEYINPUT99), .A3(new_n218_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n367_), .B(new_n368_), .C1(new_n224_), .C2(new_n211_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT104), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n356_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n371_), .B2(new_n370_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT20), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n246_), .B2(new_n356_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n353_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n370_), .A2(new_n356_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n338_), .B(new_n220_), .C1(new_n242_), .C2(new_n245_), .ZN(new_n378_));
  AND4_X1   g177(.A1(KEYINPUT20), .A2(new_n377_), .A3(new_n378_), .A4(new_n353_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n350_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n350_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n338_), .A2(new_n365_), .A3(new_n369_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n352_), .B1(new_n375_), .B2(new_n383_), .ZN(new_n384_));
  AND4_X1   g183(.A1(KEYINPUT20), .A2(new_n377_), .A3(new_n378_), .A4(new_n352_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n381_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(KEYINPUT27), .A3(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n377_), .A2(new_n378_), .A3(KEYINPUT20), .A4(new_n352_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n232_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT87), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(new_n241_), .A3(new_n229_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n338_), .B1(new_n391_), .B2(new_n220_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n392_), .A2(new_n382_), .A3(new_n374_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n388_), .B(new_n350_), .C1(new_n393_), .C2(new_n352_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n386_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n387_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n260_), .A2(new_n317_), .A3(new_n346_), .A4(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n398_), .A2(new_n316_), .A3(new_n346_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT103), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n308_), .A2(KEYINPUT33), .A3(new_n312_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n303_), .A2(new_n262_), .A3(new_n304_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n301_), .A2(new_n302_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n262_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n314_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n404_), .A2(new_n407_), .A3(KEYINPUT102), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT102), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(KEYINPUT4), .ZN(new_n410_));
  INV_X1    g209(.A(new_n304_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n306_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n312_), .B1(new_n405_), .B2(new_n262_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n403_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n314_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n386_), .B(new_n394_), .C1(new_n416_), .C2(KEYINPUT33), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n402_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n395_), .B1(new_n313_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT102), .B1(new_n404_), .B2(new_n407_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n421_), .A2(new_n422_), .B1(new_n416_), .B2(KEYINPUT33), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT103), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n384_), .A2(new_n385_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n316_), .B(new_n426_), .C1(new_n427_), .C2(new_n425_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n401_), .B1(new_n429_), .B2(new_n346_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n400_), .B1(new_n430_), .B2(new_n260_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G190gat), .B(G218gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT75), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G134gat), .B(G162gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  INV_X1    g234(.A(KEYINPUT36), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G232gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT34), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G29gat), .B(G36gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G43gat), .B(G50gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n446_), .B(new_n448_), .C1(new_n450_), .C2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT67), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  AND2_X1   g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT8), .B1(new_n453_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT65), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT65), .B1(new_n450_), .B2(new_n452_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n448_), .A2(new_n446_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n451_), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT65), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n463_), .A3(new_n467_), .A4(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT8), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n457_), .A2(new_n475_), .A3(new_n460_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n462_), .B1(new_n468_), .B2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n479_));
  INV_X1    g278(.A(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n472_), .A2(new_n473_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n454_), .B1(new_n459_), .B2(KEYINPUT9), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT64), .B1(new_n459_), .B2(KEYINPUT9), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT9), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n456_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n484_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT70), .B1(new_n483_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT70), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n484_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n466_), .A2(new_n491_), .A3(new_n492_), .A4(new_n482_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n445_), .B1(new_n478_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n461_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n475_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n474_), .A2(new_n476_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n472_), .A2(new_n467_), .A3(new_n473_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT66), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n498_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n483_), .A2(new_n489_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n502_), .A2(new_n443_), .A3(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT35), .B(new_n440_), .C1(new_n495_), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n494_), .A2(new_n478_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n445_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n440_), .A2(KEYINPUT35), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n501_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n503_), .B1(new_n510_), .B2(new_n462_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n443_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n440_), .A2(KEYINPUT35), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n508_), .A2(new_n509_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n438_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n505_), .A2(new_n515_), .A3(KEYINPUT76), .A4(new_n437_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n435_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n516_), .A2(KEYINPUT36), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(G15gat), .A2(G22gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G15gat), .A2(G22gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(G1gat), .B2(G8gat), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n526_), .A2(new_n528_), .A3(KEYINPUT78), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531_));
  INV_X1    g330(.A(G8gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT79), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT78), .B1(new_n526_), .B2(new_n528_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G1gat), .B(G8gat), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n541_), .A3(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT80), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT80), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n547_), .A3(new_n544_), .ZN(new_n548_));
  AND4_X1   g347(.A1(G231gat), .A2(new_n546_), .A3(G233gat), .A4(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT11), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  INV_X1    g352(.A(G64gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G57gat), .ZN(new_n555_));
  INV_X1    g354(.A(G57gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G64gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n546_), .A2(new_n548_), .B1(G231gat), .B2(G233gat), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n549_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n549_), .B2(new_n563_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n565_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n561_), .A2(KEYINPUT68), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n575_), .B(new_n552_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n549_), .A2(new_n577_), .A3(new_n563_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n549_), .B2(new_n563_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n570_), .B(KEYINPUT17), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n573_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n503_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n478_), .A2(new_n590_), .A3(new_n577_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n577_), .B1(new_n478_), .B2(new_n590_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT69), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n511_), .A2(KEYINPUT69), .A3(new_n577_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n589_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n562_), .A2(KEYINPUT12), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n506_), .A2(new_n598_), .B1(new_n511_), .B2(new_n577_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n511_), .B2(new_n577_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n588_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n587_), .B1(new_n596_), .B2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n602_), .A3(new_n587_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n596_), .A2(KEYINPUT71), .A3(new_n602_), .A4(new_n587_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n603_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT72), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n603_), .B(new_n613_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n545_), .A2(new_n512_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n443_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT82), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n618_), .A2(new_n619_), .A3(KEYINPUT83), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT83), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n535_), .A2(new_n541_), .A3(new_n539_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n541_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n512_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n624_), .B2(KEYINPUT82), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n617_), .B1(new_n620_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G229gat), .A2(G233gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT83), .B1(new_n618_), .B2(new_n619_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n624_), .A2(KEYINPUT82), .A3(new_n621_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n616_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(new_n628_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n545_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n618_), .B1(new_n633_), .B2(new_n507_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n627_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT84), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G169gat), .B(G197gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n638_), .B(new_n639_), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n632_), .A2(new_n635_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n615_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n431_), .A2(new_n523_), .A3(new_n582_), .A4(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n202_), .B1(new_n649_), .B2(new_n316_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n429_), .A2(new_n346_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n401_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n260_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n400_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT85), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n632_), .A2(new_n635_), .A3(new_n642_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n642_), .B1(new_n632_), .B2(new_n635_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n641_), .A2(KEYINPUT85), .A3(new_n643_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n655_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT77), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n522_), .A2(new_n663_), .A3(KEYINPUT37), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT37), .B1(new_n522_), .B2(new_n663_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n582_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT73), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT73), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n669_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n662_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT105), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n662_), .A2(new_n677_), .A3(new_n674_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n202_), .A3(new_n316_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n681_));
  AOI21_X1  g480(.A(new_n650_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n681_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n679_), .A2(new_n202_), .A3(new_n683_), .A4(new_n316_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1324gat));
  NOR2_X1   g486(.A1(new_n399_), .A2(G8gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n676_), .A2(new_n678_), .A3(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n645_), .A2(new_n399_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT39), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(G8gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n690_), .B2(G8gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT110), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n689_), .B(new_n696_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n695_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1325gat));
  NAND2_X1  g500(.A1(new_n649_), .A2(new_n260_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT41), .B1(new_n702_), .B2(G15gat), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n257_), .A2(new_n259_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(G15gat), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n703_), .A2(new_n704_), .B1(new_n675_), .B2(new_n706_), .ZN(G1326gat));
  OR3_X1    g506(.A1(new_n675_), .A2(G22gat), .A3(new_n346_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n346_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(G22gat), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G22gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n708_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT112), .ZN(G1327gat));
  NAND2_X1  g514(.A1(new_n668_), .A2(new_n522_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n615_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n662_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(G29gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n316_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n431_), .A2(new_n722_), .A3(new_n667_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n431_), .A2(KEYINPUT113), .A3(new_n722_), .A4(new_n667_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n431_), .A2(new_n667_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT43), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n644_), .A2(new_n668_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(KEYINPUT114), .A2(KEYINPUT44), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n729_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n317_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n721_), .B1(new_n735_), .B2(new_n720_), .ZN(G1328gat));
  NOR3_X1   g535(.A1(new_n718_), .A2(G36gat), .A3(new_n399_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n733_), .A2(new_n734_), .A3(new_n399_), .ZN(new_n740_));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n739_), .B(KEYINPUT46), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  INV_X1    g545(.A(G43gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n719_), .A2(new_n747_), .A3(new_n260_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n733_), .A2(new_n734_), .A3(new_n705_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n747_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT47), .B(new_n748_), .C1(new_n749_), .C2(new_n747_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1330gat));
  AOI21_X1  g553(.A(G50gat), .B1(new_n719_), .B2(new_n709_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n733_), .A2(new_n734_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n709_), .A2(G50gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(G1331gat));
  AND2_X1   g557(.A1(new_n672_), .A2(new_n673_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n582_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n655_), .A2(new_n522_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n556_), .A3(new_n317_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n641_), .A2(new_n643_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n671_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n431_), .A2(new_n669_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n316_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n764_), .B1(new_n771_), .B2(new_n556_), .ZN(G1332gat));
  OAI21_X1  g571(.A(G64gat), .B1(new_n763_), .B2(new_n399_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT48), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n554_), .A3(new_n398_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1333gat));
  OR3_X1    g575(.A1(new_n767_), .A2(G71gat), .A3(new_n705_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n761_), .A2(new_n260_), .A3(new_n762_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(G71gat), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G71gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT117), .Z(G1334gat));
  OAI21_X1  g582(.A(G78gat), .B1(new_n763_), .B2(new_n346_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n346_), .A2(G78gat), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT119), .Z(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n767_), .B2(new_n788_), .ZN(G1335gat));
  NOR3_X1   g588(.A1(new_n671_), .A2(new_n765_), .A3(new_n582_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n729_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n317_), .ZN(new_n792_));
  NOR4_X1   g591(.A1(new_n655_), .A2(new_n759_), .A3(new_n765_), .A4(new_n716_), .ZN(new_n793_));
  INV_X1    g592(.A(G85gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n316_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(G1336gat));
  OAI21_X1  g595(.A(G92gat), .B1(new_n791_), .B2(new_n399_), .ZN(new_n797_));
  INV_X1    g596(.A(G92gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n793_), .A2(new_n798_), .A3(new_n398_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n791_), .B2(new_n705_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n793_), .A2(new_n260_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n793_), .A2(new_n480_), .A3(new_n709_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n729_), .A2(new_n709_), .A3(new_n790_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(G106gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n805_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  NOR3_X1   g613(.A1(new_n398_), .A2(new_n317_), .A3(new_n709_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NOR2_X1   g615(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n588_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n602_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n599_), .A2(KEYINPUT55), .A3(new_n588_), .A4(new_n601_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n817_), .B1(new_n822_), .B2(new_n586_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n817_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n587_), .B(new_n824_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n641_), .A2(new_n643_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n608_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n626_), .A2(new_n627_), .A3(new_n631_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n642_), .B1(new_n634_), .B2(new_n628_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n643_), .A2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n826_), .A2(new_n827_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n816_), .B1(new_n833_), .B2(new_n522_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n490_), .A2(new_n493_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n598_), .B1(new_n502_), .B2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n591_), .C1(new_n592_), .C2(KEYINPUT12), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n819_), .B1(new_n837_), .B2(new_n589_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n589_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n821_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n586_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n824_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n606_), .A2(new_n607_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n822_), .A2(new_n586_), .A3(new_n817_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n843_), .A2(new_n765_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n828_), .A2(new_n832_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT57), .A3(new_n523_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n834_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n844_), .A2(new_n643_), .A3(new_n831_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n822_), .B2(new_n586_), .ZN(new_n854_));
  AOI211_X1 g653(.A(KEYINPUT56), .B(new_n587_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT58), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT121), .B1(new_n859_), .B2(KEYINPUT58), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n852_), .B2(new_n856_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n667_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n582_), .B1(new_n850_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n615_), .A2(new_n760_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n666_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n582_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n865_), .A2(new_n671_), .A3(new_n868_), .A4(new_n666_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n260_), .B(new_n815_), .C1(new_n864_), .C2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(new_n765_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n851_), .A2(new_n854_), .A3(new_n855_), .A4(KEYINPUT121), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(KEYINPUT122), .ZN(new_n879_));
  INV_X1    g678(.A(new_n862_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n666_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n834_), .A2(new_n849_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n668_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n867_), .A2(new_n869_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n885_), .A2(KEYINPUT59), .A3(new_n260_), .A4(new_n815_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n661_), .B1(new_n876_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n874_), .B1(new_n887_), .B2(new_n873_), .ZN(G1340gat));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n671_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n872_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n889_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n759_), .B1(new_n876_), .B2(new_n886_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g692(.A(G127gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n872_), .A2(new_n894_), .A3(new_n582_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n668_), .B1(new_n876_), .B2(new_n886_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(KEYINPUT123), .B(new_n895_), .C1(new_n896_), .C2(new_n894_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1342gat));
  INV_X1    g700(.A(G134gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n872_), .A2(new_n902_), .A3(new_n522_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n666_), .B1(new_n876_), .B2(new_n886_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n902_), .ZN(G1343gat));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n842_), .A2(KEYINPUT56), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n822_), .A2(new_n853_), .A3(new_n586_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(new_n832_), .A3(new_n844_), .A4(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n859_), .B1(new_n909_), .B2(KEYINPUT121), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n862_), .B1(new_n910_), .B2(new_n877_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n834_), .B(new_n849_), .C1(new_n911_), .C2(new_n666_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n870_), .B1(new_n912_), .B2(new_n668_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n705_), .A2(new_n316_), .A3(new_n709_), .A4(new_n399_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n906_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n914_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT124), .B(new_n916_), .C1(new_n864_), .C2(new_n870_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n765_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g719(.A(new_n759_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT125), .B1(new_n918_), .B2(new_n582_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927_));
  AOI211_X1 g726(.A(new_n927_), .B(new_n668_), .C1(new_n915_), .C2(new_n917_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n925_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(KEYINPUT124), .B1(new_n885_), .B2(new_n916_), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n906_), .B(new_n914_), .C1(new_n883_), .C2(new_n884_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n582_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n927_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n918_), .A2(KEYINPUT125), .A3(new_n582_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n924_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n929_), .A2(new_n935_), .ZN(G1346gat));
  INV_X1    g735(.A(new_n918_), .ZN(new_n937_));
  OAI21_X1  g736(.A(G162gat), .B1(new_n937_), .B2(new_n666_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n918_), .A2(new_n288_), .A3(new_n522_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n913_), .A2(new_n705_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n399_), .A2(new_n316_), .A3(new_n709_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n941_), .A2(new_n765_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT62), .B1(new_n943_), .B2(KEYINPUT22), .ZN(new_n944_));
  OAI21_X1  g743(.A(G169gat), .B1(new_n943_), .B2(KEYINPUT62), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n225_), .B2(new_n944_), .ZN(G1348gat));
  NAND2_X1  g746(.A1(new_n941_), .A2(new_n942_), .ZN(new_n948_));
  OAI21_X1  g747(.A(G176gat), .B1(new_n948_), .B2(new_n759_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n615_), .A2(new_n226_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(new_n950_), .ZN(G1349gat));
  OR4_X1    g750(.A1(KEYINPUT126), .A2(new_n948_), .A3(new_n243_), .A4(new_n668_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n948_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n243_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n953_), .A2(new_n954_), .A3(new_n582_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(KEYINPUT126), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n234_), .B1(new_n948_), .B2(new_n668_), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n952_), .A2(new_n956_), .A3(new_n957_), .ZN(G1350gat));
  OAI21_X1  g757(.A(G190gat), .B1(new_n948_), .B2(new_n666_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n522_), .A2(new_n233_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n948_), .B2(new_n960_), .ZN(G1351gat));
  NAND4_X1  g760(.A1(new_n705_), .A2(new_n317_), .A3(new_n709_), .A4(new_n398_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n913_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n765_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n921_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g766(.A1(new_n963_), .A2(new_n582_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(KEYINPUT63), .B(G211gat), .ZN(new_n969_));
  OR3_X1    g768(.A1(new_n968_), .A2(KEYINPUT127), .A3(new_n969_), .ZN(new_n970_));
  OAI21_X1  g769(.A(KEYINPUT127), .B1(new_n968_), .B2(new_n969_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n968_), .A2(new_n972_), .ZN(new_n973_));
  AND3_X1   g772(.A1(new_n970_), .A2(new_n971_), .A3(new_n973_), .ZN(G1354gat));
  INV_X1    g773(.A(G218gat), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n963_), .A2(new_n975_), .A3(new_n522_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n913_), .A2(new_n666_), .A3(new_n962_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n975_), .ZN(G1355gat));
endmodule


