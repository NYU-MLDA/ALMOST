//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n553_, new_n554_, new_n555_, new_n556_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n211_), .B1(new_n216_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(KEYINPUT67), .B(new_n211_), .C1(new_n216_), .C2(new_n222_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT8), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n216_), .B2(new_n222_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n213_), .A2(new_n215_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n230_), .A2(KEYINPUT65), .A3(new_n221_), .A4(new_n220_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n211_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT66), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n229_), .A2(new_n236_), .A3(new_n233_), .A4(new_n231_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT10), .B(G99gat), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n219_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(G92gat), .ZN(new_n243_));
  OR3_X1    g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT9), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n244_), .A4(new_n230_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n210_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n206_), .A2(new_n207_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n238_), .A2(new_n245_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT34), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT35), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n248_), .B1(new_n256_), .B2(KEYINPUT70), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(KEYINPUT70), .B2(new_n256_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n253_), .A2(new_n254_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n248_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n255_), .A4(new_n250_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n247_), .B1(new_n254_), .B2(new_n253_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT73), .B1(new_n263_), .B2(new_n256_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n258_), .A2(new_n259_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G190gat), .B(G218gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT71), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G134gat), .B(G162gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT36), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT36), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT72), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n265_), .A2(KEYINPUT74), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT74), .B1(new_n265_), .B2(new_n276_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT37), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT37), .B(new_n272_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G57gat), .B(G64gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT11), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT11), .ZN(new_n286_));
  XOR2_X1   g085(.A(G71gat), .B(G78gat), .Z(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT75), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n294_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n292_), .B(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G183gat), .B(G211gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT17), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(KEYINPUT76), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT17), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n302_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT76), .B1(new_n302_), .B2(new_n307_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n283_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT77), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT87), .B(G197gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(KEYINPUT21), .B(new_n319_), .C1(new_n320_), .C2(G204gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G197gat), .A2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(new_n320_), .B2(G204gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT21), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(KEYINPUT21), .ZN(new_n326_));
  OAI22_X1  g125(.A1(new_n322_), .A2(new_n325_), .B1(new_n318_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(KEYINPUT24), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT25), .B(G183gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n328_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n332_), .A2(new_n334_), .A3(new_n337_), .A4(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n334_), .B1(G183gat), .B2(G190gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT22), .B(G169gat), .Z(new_n342_));
  OAI211_X1 g141(.A(new_n341_), .B(new_n331_), .C1(G176gat), .C2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n327_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n342_), .A2(KEYINPUT83), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  INV_X1    g146(.A(G169gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT22), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n349_), .B2(KEYINPUT83), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n341_), .B(new_n331_), .C1(new_n346_), .C2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n332_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n330_), .A2(KEYINPUT24), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n345_), .B(KEYINPUT20), .C1(new_n327_), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT19), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n354_), .A2(new_n327_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n327_), .A2(new_n344_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT20), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n361_), .B2(KEYINPUT90), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(KEYINPUT90), .B2(new_n361_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n358_), .B1(new_n363_), .B2(new_n357_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT18), .ZN(new_n366_));
  XOR2_X1   g165(.A(G64gat), .B(G92gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  INV_X1    g169(.A(new_n361_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n359_), .A2(new_n357_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n371_), .A2(new_n372_), .B1(new_n357_), .B2(new_n355_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n373_), .B2(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n373_), .A2(new_n368_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n368_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n370_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G155gat), .ZN(new_n381_));
  INV_X1    g180(.A(G162gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT1), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G155gat), .A3(G162gat), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n383_), .B(new_n385_), .C1(G155gat), .C2(G162gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(G141gat), .B(G148gat), .Z(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n381_), .A2(new_n382_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT86), .ZN(new_n399_));
  AOI211_X1 g198(.A(new_n391_), .B(new_n392_), .C1(new_n397_), .C2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n390_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n327_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G78gat), .B(G106gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT89), .B1(new_n405_), .B2(new_n406_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n401_), .A2(new_n402_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G22gat), .B(G50gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT28), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n409_), .B(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n380_), .A2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G127gat), .B(G134gat), .Z(new_n418_));
  XOR2_X1   g217(.A(G113gat), .B(G120gat), .Z(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n401_), .B(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT4), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n420_), .B1(new_n390_), .B2(new_n400_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n422_), .B(new_n424_), .C1(KEYINPUT4), .C2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n421_), .A2(new_n423_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(G85gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n426_), .A2(new_n432_), .A3(new_n427_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT84), .B(G15gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n354_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(new_n420_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(G43gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT31), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n441_), .B(new_n446_), .Z(new_n447_));
  NOR2_X1   g246(.A1(new_n436_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n417_), .A2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n434_), .A2(new_n435_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n368_), .A2(KEYINPUT32), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n373_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n364_), .B2(new_n451_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n426_), .A2(KEYINPUT33), .A3(new_n432_), .A4(new_n427_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n432_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n422_), .B1(KEYINPUT4), .B2(new_n425_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n424_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n454_), .A2(new_n376_), .A3(new_n457_), .A4(new_n377_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n435_), .A2(new_n459_), .ZN(new_n460_));
  OAI22_X1  g259(.A1(new_n450_), .A2(new_n453_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n416_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n436_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n369_), .A2(new_n374_), .B1(new_n378_), .B2(new_n370_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n461_), .A2(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n447_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n449_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n238_), .A2(new_n245_), .A3(new_n290_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n290_), .B1(new_n238_), .B2(new_n245_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n473_), .B(KEYINPUT64), .Z(new_n474_));
  INV_X1    g273(.A(new_n290_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n246_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT12), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n472_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n238_), .A2(new_n245_), .A3(new_n290_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G120gat), .B(G148gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT5), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G176gat), .B(G204gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(KEYINPUT13), .A3(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT78), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n301_), .B2(new_n208_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n294_), .B(new_n299_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n249_), .A2(new_n500_), .A3(KEYINPUT78), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(new_n249_), .B2(new_n500_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n499_), .A2(new_n501_), .B1(new_n208_), .B2(new_n301_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT79), .B1(new_n508_), .B2(new_n505_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n208_), .A2(new_n209_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT15), .B1(new_n206_), .B2(new_n207_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n301_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(new_n505_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT80), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n502_), .A2(new_n512_), .A3(new_n515_), .A4(new_n505_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n507_), .A2(new_n509_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G113gat), .B(G141gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT81), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n507_), .A2(new_n509_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n514_), .A2(new_n516_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n497_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n467_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n315_), .A2(new_n529_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n530_), .A2(G1gat), .A3(new_n450_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT38), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT91), .Z(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(KEYINPUT38), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT93), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(KEYINPUT92), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n497_), .B2(new_n527_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n279_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(new_n313_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n467_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(G1gat), .B1(new_n543_), .B2(new_n450_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n533_), .A2(new_n535_), .A3(new_n544_), .ZN(G1324gat));
  AOI21_X1  g344(.A(new_n297_), .B1(new_n542_), .B2(new_n380_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT39), .Z(new_n547_));
  INV_X1    g346(.A(new_n530_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n297_), .A3(new_n380_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(KEYINPUT94), .B(KEYINPUT40), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(G1325gat));
  INV_X1    g351(.A(G15gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n542_), .B2(new_n466_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT41), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n466_), .A2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n555_), .B1(new_n530_), .B2(new_n556_), .ZN(G1326gat));
  INV_X1    g356(.A(G22gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n542_), .B2(new_n416_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT42), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n548_), .A2(new_n558_), .A3(new_n416_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT95), .Z(G1327gat));
  INV_X1    g362(.A(new_n313_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n279_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n529_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n567_), .A2(G29gat), .A3(new_n450_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT43), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n467_), .B2(new_n283_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n467_), .A2(new_n569_), .A3(new_n283_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT96), .B1(new_n539_), .B2(new_n313_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n539_), .A2(KEYINPUT96), .A3(new_n313_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n573_), .B(KEYINPUT44), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n572_), .ZN(new_n577_));
  OAI22_X1  g376(.A1(new_n577_), .A2(new_n570_), .B1(new_n575_), .B2(new_n574_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT97), .B(KEYINPUT44), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n436_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n583_), .A2(KEYINPUT98), .A3(G29gat), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT98), .B1(new_n583_), .B2(G29gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n568_), .B1(new_n584_), .B2(new_n585_), .ZN(G1328gat));
  XNOR2_X1  g385(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n587_));
  INV_X1    g386(.A(G36gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n380_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n567_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n587_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n566_), .A2(new_n588_), .A3(new_n380_), .A4(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n576_), .A2(new_n581_), .A3(new_n380_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(G36gat), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT46), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n595_), .B2(KEYINPUT46), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT100), .B(KEYINPUT46), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n595_), .A2(KEYINPUT101), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n594_), .A2(G36gat), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n590_), .A2(new_n592_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n599_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  OAI22_X1  g405(.A1(new_n597_), .A2(new_n598_), .B1(new_n600_), .B2(new_n606_), .ZN(G1329gat));
  NAND3_X1  g406(.A1(new_n582_), .A2(G43gat), .A3(new_n466_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n443_), .B1(new_n567_), .B2(new_n447_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g410(.A(G50gat), .B1(new_n566_), .B2(new_n416_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n416_), .A2(G50gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n582_), .B2(new_n613_), .ZN(G1331gat));
  INV_X1    g413(.A(new_n497_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n523_), .A2(new_n526_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n467_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n541_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT104), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n620_), .A2(G57gat), .A3(new_n436_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n315_), .A2(new_n618_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G57gat), .B1(new_n622_), .B2(new_n436_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n621_), .B1(new_n625_), .B2(new_n626_), .ZN(G1332gat));
  INV_X1    g426(.A(G64gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n620_), .B2(new_n380_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n464_), .A2(G64gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT106), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n622_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(G1333gat));
  INV_X1    g434(.A(G71gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n620_), .B2(new_n466_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT49), .Z(new_n638_));
  NOR2_X1   g437(.A1(new_n447_), .A2(G71gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT107), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n622_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(G1334gat));
  INV_X1    g441(.A(G78gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n620_), .B2(new_n416_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT50), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n622_), .A2(new_n643_), .A3(new_n416_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1335gat));
  NAND3_X1  g446(.A1(new_n573_), .A2(new_n313_), .A3(new_n617_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT109), .ZN(new_n649_));
  OAI21_X1  g448(.A(G85gat), .B1(new_n649_), .B2(new_n450_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n618_), .A2(new_n565_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT108), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n242_), .A3(new_n436_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(G1336gat));
  OAI21_X1  g453(.A(G92gat), .B1(new_n649_), .B2(new_n464_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n243_), .A3(new_n380_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1337gat));
  OAI21_X1  g456(.A(G99gat), .B1(new_n649_), .B2(new_n447_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n239_), .A3(new_n466_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT51), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT51), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n662_), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1338gat));
  NAND3_X1  g463(.A1(new_n652_), .A2(new_n219_), .A3(new_n416_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n648_), .A2(new_n462_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT52), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G106gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G106gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT53), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT53), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n672_), .B(new_n665_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1339gat));
  NAND3_X1  g473(.A1(new_n417_), .A2(new_n436_), .A3(new_n466_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT122), .Z(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT57), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n540_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n521_), .B1(new_n508_), .B2(new_n506_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n502_), .A2(new_n512_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT117), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n505_), .B1(new_n681_), .B2(KEYINPUT117), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT118), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n493_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n685_), .B2(new_n493_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n616_), .A2(new_n492_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n693_));
  NAND2_X1  g492(.A1(new_n480_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT113), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n480_), .A2(new_n696_), .A3(new_n693_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n474_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n246_), .A2(new_n475_), .B1(new_n477_), .B2(KEYINPUT12), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n482_), .B2(new_n469_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n702_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n474_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n472_), .A2(KEYINPUT55), .A3(new_n479_), .A4(new_n474_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT114), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n703_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n489_), .B1(new_n700_), .B2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n698_), .B1(new_n694_), .B2(KEYINPUT113), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n703_), .A2(new_n706_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n697_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n489_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n692_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT116), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n691_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n492_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n527_), .A2(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n489_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n709_), .B1(new_n714_), .B2(new_n489_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(KEYINPUT116), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n679_), .B1(new_n718_), .B2(new_n724_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n526_), .A2(new_n719_), .A3(new_n684_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n489_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n721_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT58), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT120), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT56), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n708_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n715_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT120), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(KEYINPUT58), .A4(new_n726_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n728_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n730_), .A2(new_n283_), .A3(new_n735_), .A4(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n690_), .B1(new_n723_), .B2(KEYINPUT116), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n716_), .A2(new_n717_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n540_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n725_), .B(new_n738_), .C1(new_n741_), .C2(KEYINPUT57), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT121), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n279_), .B1(new_n718_), .B2(new_n724_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n678_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n746_), .A2(KEYINPUT121), .A3(new_n725_), .A4(new_n738_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n747_), .A3(new_n313_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n495_), .A2(new_n527_), .A3(new_n564_), .A4(new_n496_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(KEYINPUT110), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(KEYINPUT110), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n752_), .B(new_n283_), .C1(KEYINPUT111), .C2(KEYINPUT54), .ZN(new_n753_));
  INV_X1    g552(.A(new_n283_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n752_), .ZN(new_n755_));
  OR2_X1    g554(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n756_));
  NAND2_X1  g555(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n754_), .A2(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n753_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n677_), .B1(new_n748_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n616_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n753_), .A2(new_n758_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n564_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n747_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT59), .B1(new_n765_), .B2(new_n677_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n742_), .A2(new_n313_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n759_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n677_), .A2(KEYINPUT59), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n766_), .A2(new_n616_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n762_), .B1(new_n772_), .B2(new_n761_), .ZN(G1340gat));
  INV_X1    g572(.A(KEYINPUT124), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT123), .ZN(new_n775_));
  AND2_X1   g574(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n776_));
  NOR2_X1   g575(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n497_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n760_), .B2(new_n779_), .ZN(new_n780_));
  NOR4_X1   g579(.A1(new_n765_), .A2(KEYINPUT123), .A3(new_n677_), .A4(new_n778_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(G120gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n615_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n766_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n774_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n748_), .A2(new_n759_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n676_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n770_), .A2(new_n497_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G120gat), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(KEYINPUT124), .C1(new_n780_), .C2(new_n781_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n786_), .A2(new_n792_), .ZN(G1341gat));
  INV_X1    g592(.A(G127gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n760_), .A2(new_n794_), .A3(new_n564_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n766_), .A2(new_n564_), .A3(new_n770_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n794_), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n760_), .A2(new_n799_), .A3(new_n540_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n766_), .A2(new_n283_), .A3(new_n770_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(new_n799_), .ZN(G1343gat));
  NOR4_X1   g602(.A1(new_n462_), .A2(new_n380_), .A3(new_n450_), .A4(new_n466_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n788_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n616_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n497_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g609(.A(KEYINPUT61), .B(G155gat), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT125), .B1(new_n805_), .B2(new_n313_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n805_), .A2(KEYINPUT125), .A3(new_n313_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OR3_X1    g615(.A1(new_n805_), .A2(KEYINPUT125), .A3(new_n313_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n813_), .A3(new_n811_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1346gat));
  OAI21_X1  g618(.A(G162gat), .B1(new_n805_), .B2(new_n754_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n540_), .A2(new_n382_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n805_), .B2(new_n821_), .ZN(G1347gat));
  AOI21_X1  g621(.A(new_n416_), .B1(new_n759_), .B2(new_n767_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n380_), .A2(new_n448_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(G169gat), .B1(new_n826_), .B2(new_n527_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n828_), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n826_), .A2(new_n342_), .A3(new_n527_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(G1348gat));
  NOR2_X1   g631(.A1(new_n765_), .A2(new_n416_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n824_), .A2(new_n347_), .A3(new_n615_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n823_), .A2(new_n497_), .A3(new_n825_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n833_), .A2(new_n834_), .B1(new_n835_), .B2(new_n347_), .ZN(G1349gat));
  NOR2_X1   g635(.A1(new_n824_), .A2(new_n313_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G183gat), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n824_), .A2(new_n313_), .A3(new_n335_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n823_), .B2(new_n839_), .ZN(G1350gat));
  NAND4_X1  g639(.A1(new_n823_), .A2(new_n540_), .A3(new_n336_), .A4(new_n825_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n826_), .A2(new_n754_), .ZN(new_n842_));
  INV_X1    g641(.A(G190gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT126), .B(new_n841_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1351gat));
  AND3_X1   g647(.A1(new_n463_), .A2(new_n380_), .A3(new_n447_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n788_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(G197gat), .A3(new_n616_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT127), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(G197gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n788_), .A2(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n527_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n850_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n616_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n853_), .A2(new_n856_), .A3(new_n857_), .ZN(G1352gat));
  NAND2_X1  g657(.A1(new_n850_), .A2(new_n497_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  AND2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n855_), .A2(new_n313_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n850_), .A2(new_n564_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n861_), .ZN(G1354gat));
  OR3_X1    g664(.A1(new_n855_), .A2(G218gat), .A3(new_n279_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G218gat), .B1(new_n855_), .B2(new_n754_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1355gat));
endmodule


