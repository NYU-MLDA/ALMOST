//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT69), .B(G71gat), .ZN(new_n205_));
  INV_X1    g004(.A(G78gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n204_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT69), .B(G71gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G78gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(KEYINPUT11), .A3(new_n207_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G57gat), .B(G64gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n214_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(KEYINPUT11), .A3(new_n207_), .A4(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n220_));
  OAI22_X1  g019(.A1(new_n219_), .A2(new_n220_), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n221_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G85gat), .B(G92gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n231_), .A2(new_n238_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT10), .B(G99gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT9), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n242_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT9), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n243_), .A2(new_n248_), .ZN(new_n250_));
  NOR4_X1   g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT65), .A4(new_n245_), .ZN(new_n251_));
  OAI221_X1 g050(.A(new_n226_), .B1(G106gat), .B2(new_n241_), .C1(new_n247_), .C2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n218_), .B1(new_n240_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n253_), .B2(KEYINPUT12), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n240_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n218_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT71), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n255_), .A2(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n240_), .A2(KEYINPUT70), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n235_), .A2(new_n237_), .A3(new_n263_), .A4(new_n239_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n252_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n218_), .A2(new_n258_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n261_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n260_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n261_), .B2(new_n253_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G120gat), .B(G148gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT5), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G176gat), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n273_), .A2(new_n278_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n202_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n279_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT72), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G15gat), .B(G22gat), .ZN(new_n287_));
  INV_X1    g086(.A(G1gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n218_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT80), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT16), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(G183gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G211gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(KEYINPUT17), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n296_), .B1(KEYINPUT79), .B2(new_n302_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(KEYINPUT79), .B2(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G29gat), .B(G36gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(G43gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(G43gat), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(G50gat), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(G50gat), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT74), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n310_), .ZN(new_n314_));
  INV_X1    g113(.A(G50gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(G50gat), .A3(new_n310_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n313_), .A2(new_n319_), .A3(KEYINPUT15), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT15), .B1(new_n313_), .B2(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n252_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n316_), .A2(new_n317_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT76), .B1(new_n255_), .B2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G232gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT34), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n330_), .A2(new_n331_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n330_), .B(new_n331_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G190gat), .B(G218gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT75), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(G134gat), .ZN(new_n339_));
  INV_X1    g138(.A(G162gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT36), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(KEYINPUT36), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n336_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n336_), .A2(new_n343_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n336_), .A2(KEYINPUT77), .A3(new_n343_), .A4(new_n344_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n345_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT37), .B1(new_n353_), .B2(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n286_), .A2(new_n307_), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G113gat), .B(G141gat), .ZN(new_n358_));
  INV_X1    g157(.A(G169gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G197gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n326_), .A2(new_n293_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G229gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT81), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n320_), .A2(new_n321_), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n363_), .B(new_n365_), .C1(new_n366_), .C2(new_n293_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n326_), .B(new_n293_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(G229gat), .A3(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n362_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n363_), .B1(new_n366_), .B2(new_n293_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n365_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n362_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n376_), .A3(KEYINPUT82), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT82), .B1(new_n371_), .B2(new_n376_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OR2_X1    g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  INV_X1    g181(.A(G141gat), .ZN(new_n383_));
  INV_X1    g182(.A(G148gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n385_), .A2(KEYINPUT3), .B1(new_n386_), .B2(KEYINPUT92), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT89), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(G141gat), .A3(G148gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT2), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n386_), .A2(KEYINPUT92), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n385_), .A2(KEYINPUT3), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n381_), .B(new_n382_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n398_));
  OR3_X1    g197(.A1(new_n382_), .A2(new_n398_), .A3(KEYINPUT1), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n382_), .B2(KEYINPUT1), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n382_), .A2(KEYINPUT1), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(new_n381_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n385_), .B(KEYINPUT90), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n402_), .A2(new_n389_), .A3(new_n403_), .A4(new_n391_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G127gat), .ZN(new_n406_));
  INV_X1    g205(.A(G134gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G127gat), .A2(G134gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n413_));
  OAI21_X1  g212(.A(G113gat), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT88), .ZN(new_n416_));
  INV_X1    g215(.A(G113gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n411_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(G120gat), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(G120gat), .B1(new_n414_), .B2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n405_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(G120gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(new_n404_), .A3(new_n419_), .A4(new_n397_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n426_), .A3(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n405_), .B(new_n430_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n429_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n422_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G85gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G1gat), .B(G29gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT102), .B(G57gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n434_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n432_), .A2(new_n442_), .A3(new_n433_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G183gat), .A2(G190gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT83), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G183gat), .A3(G190gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT23), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(KEYINPUT23), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT84), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n459_), .B(new_n456_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT25), .B(G183gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT26), .B(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G176gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n359_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G169gat), .A2(G176gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT24), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n458_), .A2(new_n460_), .A3(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(G183gat), .A2(G190gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n448_), .A2(new_n452_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n449_), .A2(new_n451_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n470_), .B(new_n471_), .C1(new_n472_), .C2(new_n452_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G169gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n469_), .A2(KEYINPUT85), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n455_), .A2(new_n457_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n459_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n468_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n455_), .A2(KEYINPUT84), .A3(new_n457_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n479_), .B1(new_n484_), .B2(new_n476_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n447_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT85), .B1(new_n469_), .B2(new_n477_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n479_), .A3(new_n476_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT30), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n446_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT86), .B(G43gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(G15gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n493_), .B(new_n496_), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT31), .B1(new_n490_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n487_), .A2(KEYINPUT30), .A3(new_n488_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT30), .B1(new_n487_), .B2(new_n488_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT87), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n497_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n420_), .A2(new_n421_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n499_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n486_), .A2(new_n446_), .A3(new_n489_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n490_), .A2(KEYINPUT31), .A3(new_n498_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n503_), .B1(new_n502_), .B2(new_n497_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n505_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n499_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n445_), .B1(new_n510_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT21), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n361_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(G197gat), .B2(new_n277_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n277_), .A2(G197gat), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n518_), .B(new_n519_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n361_), .A2(G204gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n361_), .A2(G204gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(new_n520_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n528_), .A2(KEYINPUT94), .A3(new_n518_), .A4(new_n519_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G211gat), .B(G218gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT21), .B1(new_n522_), .B2(new_n527_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n528_), .A2(new_n519_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n518_), .B1(new_n536_), .B2(KEYINPUT96), .ZN(new_n537_));
  INV_X1    g336(.A(new_n531_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n537_), .B(new_n538_), .C1(KEYINPUT96), .C2(new_n536_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n530_), .A2(KEYINPUT95), .A3(new_n531_), .A4(new_n532_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n405_), .A2(KEYINPUT29), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(G228gat), .A3(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(G228gat), .ZN(new_n545_));
  INV_X1    g344(.A(G233gat), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n541_), .B(new_n542_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G78gat), .B(G106gat), .Z(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n405_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n405_), .B2(KEYINPUT29), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G22gat), .B(G50gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n544_), .A2(new_n547_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n548_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n549_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n560_), .A2(new_n549_), .A3(new_n556_), .A4(KEYINPUT97), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G8gat), .B(G36gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT18), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G64gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(G92gat), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n484_), .A2(new_n476_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n541_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G226gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT19), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n475_), .B(KEYINPUT99), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n455_), .A2(new_n470_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n471_), .B1(new_n472_), .B2(new_n452_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n468_), .A2(new_n577_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n575_), .A2(new_n576_), .B1(new_n457_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n579_), .A2(new_n535_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n580_));
  AND4_X1   g379(.A1(KEYINPUT20), .A2(new_n571_), .A3(new_n574_), .A4(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n573_), .B(KEYINPUT98), .Z(new_n582_));
  INV_X1    g381(.A(KEYINPUT20), .ZN(new_n583_));
  INV_X1    g382(.A(new_n579_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n541_), .B2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n469_), .A2(new_n477_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n586_), .A2(new_n535_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n582_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n569_), .B1(new_n581_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n541_), .A2(new_n584_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(KEYINPUT20), .A3(new_n587_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n583_), .B1(new_n541_), .B2(new_n570_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n568_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n589_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT27), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n591_), .A2(new_n592_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n574_), .B1(new_n594_), .B2(new_n580_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n569_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(KEYINPUT27), .A3(new_n596_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n564_), .A2(new_n599_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT103), .B1(new_n517_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n563_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n551_), .A2(new_n556_), .B1(new_n560_), .B2(new_n549_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n599_), .A2(new_n603_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n509_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n514_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n610_), .A2(new_n611_), .A3(new_n614_), .A4(new_n445_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n589_), .A2(new_n596_), .A3(KEYINPUT100), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT100), .B1(new_n589_), .B2(new_n596_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n427_), .A2(new_n428_), .A3(new_n431_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n422_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n440_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT33), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n443_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n432_), .A2(KEYINPUT33), .A3(new_n442_), .A4(new_n433_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n616_), .A2(new_n617_), .A3(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT32), .B(new_n568_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n568_), .A2(KEYINPUT32), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n593_), .A2(new_n627_), .A3(new_n595_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n444_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n564_), .B1(new_n625_), .B2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n599_), .A2(new_n603_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n445_), .A3(new_n608_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n614_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n605_), .A2(new_n615_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n357_), .A2(new_n380_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT104), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n288_), .A3(new_n444_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT105), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n347_), .A2(new_n350_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n349_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n307_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n637_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n380_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT106), .B1(new_n649_), .B2(new_n285_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n285_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n648_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n288_), .B1(new_n654_), .B2(new_n444_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n640_), .B1(new_n641_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n643_), .A2(new_n656_), .ZN(G1324gat));
  AOI21_X1  g456(.A(new_n289_), .B1(new_n654_), .B2(new_n609_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n632_), .A2(G8gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n639_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT40), .ZN(G1325gat));
  AOI21_X1  g462(.A(new_n495_), .B1(new_n654_), .B2(new_n614_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n614_), .A2(new_n495_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n638_), .B2(new_n666_), .ZN(G1326gat));
  INV_X1    g466(.A(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n654_), .B2(new_n608_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n608_), .A2(new_n668_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n638_), .B2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(new_n307_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n645_), .A2(new_n674_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n637_), .A2(new_n651_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(G29gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n677_), .A3(new_n444_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n605_), .A2(new_n615_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n617_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n589_), .A2(new_n596_), .A3(KEYINPUT100), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n680_), .A2(new_n623_), .A3(new_n622_), .A4(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n608_), .B1(new_n682_), .B2(new_n629_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n609_), .A2(new_n564_), .A3(new_n444_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n635_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n355_), .B1(new_n679_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT110), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  INV_X1    g490(.A(new_n687_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(new_n692_), .C1(new_n636_), .C2(new_n355_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n690_), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n674_), .B1(new_n653_), .B2(new_n650_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n696_), .B2(KEYINPUT111), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n699_), .B(new_n700_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n445_), .B1(new_n698_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n678_), .B1(new_n703_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n676_), .A2(new_n705_), .A3(new_n609_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT45), .Z(new_n707_));
  OAI21_X1  g506(.A(new_n609_), .B1(new_n697_), .B2(new_n701_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n711_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n709_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1329gat));
  OAI21_X1  g515(.A(new_n614_), .B1(new_n697_), .B2(new_n701_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n635_), .A2(G43gat), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n717_), .A2(G43gat), .B1(new_n676_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g519(.A1(new_n676_), .A2(new_n315_), .A3(new_n608_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n564_), .B1(new_n698_), .B2(new_n702_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n315_), .ZN(G1331gat));
  NOR2_X1   g522(.A1(new_n636_), .A2(new_n380_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n647_), .A3(new_n286_), .ZN(new_n725_));
  INV_X1    g524(.A(G57gat), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n445_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n724_), .B(KEYINPUT113), .ZN(new_n728_));
  AND4_X1   g527(.A1(new_n285_), .A2(new_n728_), .A3(new_n674_), .A4(new_n355_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n444_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n727_), .B1(new_n730_), .B2(new_n726_), .ZN(G1332gat));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n729_), .A2(new_n732_), .A3(new_n609_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G64gat), .B1(new_n725_), .B2(new_n632_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n725_), .B2(new_n635_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT114), .Z(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n729_), .A2(new_n740_), .A3(new_n614_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1334gat));
  NAND3_X1  g541(.A1(new_n729_), .A2(new_n206_), .A3(new_n608_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G78gat), .B1(new_n725_), .B2(new_n564_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT50), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1335gat));
  AND3_X1   g545(.A1(new_n728_), .A2(new_n286_), .A3(new_n675_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n444_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n285_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n674_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n694_), .A2(new_n649_), .A3(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n444_), .A2(G85gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n747_), .B2(new_n609_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n609_), .A2(G92gat), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT115), .Z(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n751_), .B2(new_n756_), .ZN(G1337gat));
  AOI21_X1  g556(.A(new_n228_), .B1(new_n751_), .B2(new_n614_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n635_), .A2(new_n241_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n747_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g560(.A1(new_n747_), .A2(new_n229_), .A3(new_n608_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n694_), .A2(new_n649_), .A3(new_n608_), .A4(new_n750_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n254_), .A2(new_n259_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n267_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n324_), .A2(new_n772_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n271_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT118), .B(new_n271_), .C1(new_n771_), .C2(new_n773_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n270_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n260_), .A2(new_n268_), .A3(KEYINPUT55), .A4(new_n269_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n776_), .A2(new_n777_), .A3(new_n779_), .A4(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n278_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n278_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n781_), .A2(new_n278_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(KEYINPUT121), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n375_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT120), .Z(new_n791_));
  NAND2_X1  g590(.A1(new_n372_), .A2(new_n365_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n376_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n283_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n789_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n770_), .B1(new_n786_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n785_), .B2(KEYINPUT121), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(KEYINPUT58), .C1(new_n785_), .C2(new_n784_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n356_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT122), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  INV_X1    g603(.A(new_n379_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n377_), .A3(new_n283_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n785_), .B2(KEYINPUT119), .ZN(new_n807_));
  INV_X1    g606(.A(new_n785_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n782_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n283_), .A2(new_n279_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n807_), .A2(new_n810_), .B1(new_n811_), .B2(new_n794_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n804_), .B1(new_n812_), .B2(new_n646_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n807_), .A2(new_n810_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n811_), .A2(new_n794_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n645_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n798_), .A2(KEYINPUT122), .A3(new_n800_), .A4(new_n356_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n803_), .A2(new_n813_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n307_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n355_), .A2(new_n649_), .A3(new_n749_), .A4(new_n674_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(KEYINPUT54), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n307_), .B(new_n380_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(KEYINPUT117), .A3(new_n824_), .A4(new_n749_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(KEYINPUT54), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n822_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT123), .B1(new_n819_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n827_), .C1(new_n818_), .C2(new_n307_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n635_), .A2(new_n445_), .A3(new_n604_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834_), .B2(new_n380_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n816_), .A2(new_n813_), .A3(new_n801_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n828_), .B1(new_n836_), .B2(new_n674_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n829_), .A2(new_n831_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n832_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n842_), .B2(KEYINPUT59), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n649_), .A2(new_n417_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n835_), .B1(new_n843_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n286_), .B(new_n839_), .C1(new_n834_), .C2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT60), .B1(new_n285_), .B2(new_n424_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .A4(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G120gat), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1341gat));
  AOI21_X1  g652(.A(G127gat), .B1(new_n834_), .B2(new_n674_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n406_), .B1(new_n674_), .B2(new_n855_), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n840_), .B(new_n856_), .C1(new_n842_), .C2(KEYINPUT59), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n406_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n834_), .B2(new_n646_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n355_), .A2(new_n407_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n843_), .B2(new_n861_), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n609_), .A2(new_n564_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n841_), .A2(new_n444_), .A3(new_n635_), .A4(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n383_), .A3(new_n380_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G141gat), .B1(new_n864_), .B2(new_n649_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n384_), .A3(new_n286_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n286_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G148gat), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1345gat));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n864_), .B2(new_n307_), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n829_), .A2(new_n831_), .A3(new_n445_), .A4(new_n614_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n876_), .A2(new_n674_), .A3(new_n863_), .A4(new_n873_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1346gat));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n646_), .A3(new_n863_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n355_), .A2(new_n340_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n879_), .A2(new_n340_), .B1(new_n865_), .B2(new_n880_), .ZN(G1347gat));
  NOR3_X1   g680(.A1(new_n517_), .A2(new_n608_), .A3(new_n632_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n837_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n380_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G169gat), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n883_), .A2(KEYINPUT22), .A3(new_n649_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n885_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n359_), .B2(new_n889_), .ZN(G1348gat));
  INV_X1    g690(.A(new_n882_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n829_), .A2(new_n831_), .A3(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(G176gat), .A3(new_n286_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n464_), .B1(new_n883_), .B2(new_n749_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n893_), .A2(new_n897_), .A3(G176gat), .A4(new_n286_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n895_), .A2(new_n896_), .A3(new_n898_), .ZN(G1349gat));
  AOI21_X1  g698(.A(G183gat), .B1(new_n893_), .B2(new_n674_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n883_), .A2(new_n307_), .A3(new_n461_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n883_), .B2(new_n355_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n646_), .A2(new_n462_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n883_), .B2(new_n904_), .ZN(G1351gat));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n632_), .A2(new_n444_), .A3(new_n564_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n841_), .A2(new_n380_), .A3(new_n635_), .A4(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n908_), .B2(new_n361_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n361_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n907_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n829_), .A2(new_n831_), .A3(new_n614_), .A4(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n912_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n380_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n909_), .A2(new_n910_), .A3(new_n913_), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n286_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g715(.A(new_n307_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT127), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n912_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921_));
  INV_X1    g720(.A(G211gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n920_), .B(new_n923_), .ZN(G1354gat));
  AOI21_X1  g723(.A(G218gat), .B1(new_n912_), .B2(new_n646_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n356_), .A2(G218gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n912_), .B2(new_n926_), .ZN(G1355gat));
endmodule


