//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT84), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n218_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT22), .B1(new_n218_), .B2(KEYINPUT83), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n212_), .A2(new_n223_), .A3(new_n214_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n216_), .A2(new_n217_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n208_), .A2(new_n226_), .A3(KEYINPUT23), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n208_), .B2(KEYINPUT23), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n211_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT25), .B(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT81), .ZN(new_n232_));
  INV_X1    g031(.A(G190gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(KEYINPUT26), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(KEYINPUT26), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n231_), .A2(new_n234_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n218_), .A2(new_n220_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT24), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n230_), .A2(new_n238_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n225_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT85), .Z(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT30), .B(G99gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(KEYINPUT85), .ZN(new_n247_));
  INV_X1    g046(.A(new_n245_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G15gat), .B(G43gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT31), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(G71gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(new_n249_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n207_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n206_), .A3(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT90), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT86), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(G141gat), .A3(G148gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT2), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n265_), .A2(new_n270_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n271_), .A2(new_n274_), .A3(new_n276_), .A4(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G155gat), .ZN(new_n279_));
  INV_X1    g078(.A(G162gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n272_), .B1(new_n286_), .B2(KEYINPUT1), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n281_), .A2(new_n288_), .A3(new_n282_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n269_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT87), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT87), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n269_), .A2(new_n287_), .A3(new_n289_), .A4(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n285_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT29), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G228gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G211gat), .B(G218gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT21), .ZN(new_n300_));
  OR3_X1    g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G204gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(G197gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(G197gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT21), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n300_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n299_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT89), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n297_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n296_), .A2(new_n311_), .A3(new_n308_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n308_), .A2(KEYINPUT89), .B1(G228gat), .B2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(new_n285_), .B2(new_n294_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n315_), .B2(new_n309_), .ZN(new_n316_));
  AOI211_X1 g115(.A(new_n261_), .B(new_n264_), .C1(new_n312_), .C2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n311_), .B1(new_n296_), .B2(new_n308_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n315_), .A2(new_n313_), .A3(new_n309_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n263_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n316_), .A3(new_n264_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G22gat), .B(G50gat), .Z(new_n325_));
  NOR3_X1   g124(.A1(new_n295_), .A2(KEYINPUT29), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n284_), .A2(new_n278_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(new_n314_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n324_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n325_), .B1(new_n295_), .B2(KEYINPUT29), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n314_), .A3(new_n327_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n323_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n317_), .B1(new_n322_), .B2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n330_), .A2(new_n333_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(new_n261_), .A3(new_n321_), .A4(new_n320_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G92gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT18), .B(G64gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT32), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT19), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n348_));
  INV_X1    g147(.A(new_n211_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n209_), .A2(KEYINPUT82), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n227_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n348_), .B1(new_n351_), .B2(new_n213_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n230_), .A2(KEYINPUT95), .A3(new_n214_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n217_), .B(KEYINPUT93), .ZN(new_n354_));
  OR2_X1    g153(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n355_), .A2(KEYINPUT94), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT94), .B1(new_n355_), .B2(new_n356_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n220_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n231_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n241_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT92), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(KEYINPUT92), .A3(new_n241_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n240_), .A3(new_n212_), .A4(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n367_), .A3(new_n309_), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT103), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n243_), .A2(new_n308_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n368_), .A2(KEYINPUT103), .A3(new_n369_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n347_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n309_), .B1(new_n360_), .B2(new_n367_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n243_), .A2(new_n308_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n347_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n344_), .B1(new_n376_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n360_), .A2(new_n367_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n379_), .B1(new_n384_), .B2(new_n308_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n378_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n347_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n368_), .A2(new_n371_), .A3(KEYINPUT20), .A4(new_n347_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT101), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n344_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n344_), .A2(new_n391_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G1gat), .B(G29gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT99), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G57gat), .B(G85gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n285_), .A2(new_n294_), .A3(new_n204_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT96), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n204_), .B1(new_n285_), .B2(new_n294_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  INV_X1    g205(.A(new_n204_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n295_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT4), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n291_), .A2(new_n293_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT2), .B1(new_n266_), .B2(new_n268_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n277_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n413_), .A2(new_n275_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n283_), .B1(new_n415_), .B2(new_n274_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n407_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT97), .B1(new_n417_), .B2(KEYINPUT4), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT97), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n404_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n411_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n410_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n411_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n401_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n411_), .ZN(new_n426_));
  NOR4_X1   g225(.A1(new_n328_), .A2(KEYINPUT97), .A3(KEYINPUT4), .A4(new_n204_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n419_), .B1(new_n404_), .B2(new_n420_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n417_), .A2(KEYINPUT96), .A3(new_n402_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n420_), .B1(new_n430_), .B2(new_n408_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n424_), .B(new_n401_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n383_), .B(new_n394_), .C1(new_n425_), .C2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n342_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n388_), .B(new_n343_), .C1(new_n380_), .C2(new_n347_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n426_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n398_), .B(new_n399_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT100), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT100), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n411_), .B1(new_n430_), .B2(new_n408_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n401_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n426_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n410_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n423_), .A2(KEYINPUT33), .A3(new_n424_), .A4(new_n401_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n437_), .A2(new_n439_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n338_), .B1(new_n434_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n424_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n441_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n335_), .A2(new_n453_), .A3(new_n432_), .A4(new_n337_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n436_), .A2(KEYINPUT27), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n374_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n381_), .B1(new_n456_), .B2(new_n347_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n457_), .B2(new_n342_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT27), .B1(new_n435_), .B2(new_n436_), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n454_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n260_), .B1(new_n451_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n453_), .A2(new_n432_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n260_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n338_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n458_), .A2(new_n459_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G29gat), .B(G36gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G43gat), .B(G50gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G29gat), .B(G36gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT79), .B1(new_n475_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT15), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n474_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n482_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n480_), .A2(new_n481_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n480_), .A2(new_n481_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n470_), .A4(new_n473_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n488_), .A3(new_n489_), .A4(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n482_), .A2(new_n474_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n489_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n482_), .A2(KEYINPUT77), .A3(new_n474_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n496_), .A2(KEYINPUT78), .A3(new_n497_), .A4(new_n498_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n493_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G169gat), .B(G197gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n493_), .A2(new_n501_), .A3(new_n502_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n507_), .A2(KEYINPUT80), .A3(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(G99gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT10), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G99gat), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n517_), .A2(new_n519_), .A3(KEYINPUT64), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT64), .B1(new_n517_), .B2(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n515_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT6), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT66), .B(G92gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n525_), .A3(G92gat), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n522_), .A2(new_n524_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n531_));
  OR4_X1    g330(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n516_), .A3(new_n515_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT7), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n524_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n537_));
  XOR2_X1   g336(.A(G85gat), .B(G92gat), .Z(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n531_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n542_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n541_), .A2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n548_), .B(new_n531_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(KEYINPUT12), .A3(new_n551_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n541_), .A2(new_n557_), .A3(new_n549_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n553_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT5), .B(G176gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n555_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n553_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n564_), .B1(new_n554_), .B2(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n566_), .A2(new_n569_), .A3(KEYINPUT69), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT69), .B1(new_n566_), .B2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT13), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n514_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n467_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n541_), .A2(new_n474_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT35), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n541_), .A2(new_n486_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n578_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n581_), .A2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT72), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT73), .ZN(new_n594_));
  INV_X1    g393(.A(new_n586_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n578_), .A2(new_n595_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n587_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n590_), .B(KEYINPUT36), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n587_), .B2(new_n596_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT74), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(KEYINPUT74), .A3(KEYINPUT37), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n548_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n482_), .B(KEYINPUT75), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G211gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT16), .B(G183gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(KEYINPUT17), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n610_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(KEYINPUT76), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n610_), .A2(new_n615_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(KEYINPUT76), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n606_), .A2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n577_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n477_), .A3(new_n462_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT104), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT38), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n576_), .A2(new_n621_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n601_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(new_n467_), .A3(new_n631_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n462_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n627_), .A2(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(new_n465_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n624_), .A2(new_n478_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n633_), .B2(new_n465_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n642_), .B(new_n644_), .ZN(G1325gat));
  INV_X1    g444(.A(G15gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n260_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n624_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n633_), .A2(new_n260_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT41), .B1(new_n649_), .B2(G15gat), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT41), .B(G15gat), .C1(new_n633_), .C2(new_n260_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT107), .ZN(G1326gat));
  OAI21_X1  g453(.A(G22gat), .B1(new_n633_), .B2(new_n464_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT42), .ZN(new_n656_));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n624_), .A2(new_n657_), .A3(new_n338_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1327gat));
  NOR2_X1   g458(.A1(new_n621_), .A2(new_n632_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n577_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(G29gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n462_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT110), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n665_));
  INV_X1    g464(.A(new_n605_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT37), .B1(new_n601_), .B2(KEYINPUT74), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n461_), .B2(new_n466_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n621_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n671_), .A2(new_n576_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n670_), .B1(new_n467_), .B2(new_n606_), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT43), .B(new_n668_), .C1(new_n461_), .C2(new_n466_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n576_), .B(new_n676_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n674_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n665_), .B1(new_n682_), .B2(new_n462_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT109), .B(new_n634_), .C1(new_n677_), .C2(new_n681_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n664_), .B1(new_n685_), .B2(G29gat), .ZN(new_n686_));
  NOR4_X1   g485(.A1(new_n683_), .A2(new_n684_), .A3(KEYINPUT110), .A4(new_n662_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n663_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n682_), .B2(new_n637_), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT111), .B(new_n465_), .C1(new_n677_), .C2(new_n681_), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n637_), .A2(KEYINPUT112), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n637_), .A2(KEYINPUT112), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n661_), .A2(new_n693_), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  OAI21_X1  g499(.A(new_n689_), .B1(new_n694_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n691_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n682_), .A2(new_n690_), .A3(new_n637_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(G36gat), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n700_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(KEYINPUT46), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1329gat));
  INV_X1    g506(.A(G43gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n661_), .A2(new_n708_), .A3(new_n647_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n260_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(new_n708_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g511(.A(G50gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n661_), .A2(new_n713_), .A3(new_n338_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n464_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n713_), .ZN(G1331gat));
  NAND2_X1  g515(.A1(new_n573_), .A2(new_n575_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n513_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT80), .B1(new_n507_), .B2(new_n509_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(new_n467_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n621_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n668_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n462_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n723_), .A2(new_n632_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n462_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(G57gat), .B2(new_n727_), .ZN(G1332gat));
  INV_X1    g527(.A(G64gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n729_), .A3(new_n698_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n723_), .A2(new_n632_), .A3(new_n698_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n731_), .B2(G64gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n724_), .A2(new_n737_), .A3(new_n647_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n726_), .B2(new_n647_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT49), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n739_), .A2(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1334gat));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n724_), .A2(new_n744_), .A3(new_n338_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n726_), .A2(new_n338_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(G78gat), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT50), .B(new_n744_), .C1(new_n726_), .C2(new_n338_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1335gat));
  AND2_X1   g549(.A1(new_n722_), .A2(new_n660_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n462_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n671_), .A2(new_n622_), .A3(new_n721_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n634_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n754_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n751_), .B2(new_n637_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n753_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n698_), .A2(new_n527_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n753_), .B2(new_n260_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n751_), .B(new_n647_), .C1(new_n521_), .C2(new_n520_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n751_), .A2(new_n515_), .A3(new_n338_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n757_), .A2(new_n338_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G106gat), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n765_), .B(G106gat), .C1(new_n753_), .C2(new_n464_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n764_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  NAND4_X1  g573(.A1(new_n647_), .A2(new_n465_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n560_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n556_), .A2(new_n567_), .A3(new_n558_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n568_), .A2(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n564_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT114), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n566_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n514_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n781_), .A2(new_n786_), .A3(new_n564_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n484_), .A2(new_n488_), .A3(new_n497_), .A4(new_n492_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n496_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n506_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n509_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n785_), .A2(new_n790_), .B1(new_n572_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n776_), .B1(new_n796_), .B2(new_n601_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n572_), .A2(new_n795_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n784_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n720_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n787_), .B2(KEYINPUT115), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n804_));
  NOR2_X1   g603(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n782_), .A2(new_n804_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n781_), .A2(new_n564_), .A3(new_n805_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n807_), .A2(new_n566_), .A3(new_n795_), .A4(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n808_), .A2(new_n566_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(KEYINPUT58), .A3(new_n795_), .A4(new_n807_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n606_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n797_), .A2(new_n803_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT117), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n797_), .A2(new_n817_), .A3(new_n803_), .A4(new_n814_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n816_), .A2(new_n622_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n623_), .A2(new_n514_), .A3(new_n717_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT54), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n775_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n720_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n815_), .A2(new_n622_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(new_n821_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n826_), .A2(KEYINPUT59), .A3(new_n775_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT118), .B1(new_n822_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  INV_X1    g629(.A(new_n821_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n818_), .A2(new_n622_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n816_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n830_), .B(KEYINPUT59), .C1(new_n833_), .C2(new_n775_), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n824_), .B(new_n827_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n823_), .B1(new_n835_), .B2(new_n720_), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n717_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n822_), .B(new_n838_), .C1(KEYINPUT60), .C2(new_n837_), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n717_), .B(new_n827_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n837_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n822_), .B2(new_n621_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n622_), .B(new_n827_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g643(.A(G134gat), .B1(new_n822_), .B2(new_n601_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n668_), .B(new_n827_), .C1(new_n829_), .C2(new_n834_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G134gat), .ZN(G1343gat));
  AOI211_X1 g646(.A(new_n464_), .B(new_n647_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n698_), .A2(new_n634_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n720_), .A4(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n802_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n802_), .B2(new_n632_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n817_), .B1(new_n854_), .B2(new_n814_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n818_), .A2(new_n622_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n821_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(new_n338_), .A3(new_n260_), .A4(new_n850_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT120), .B1(new_n858_), .B2(new_n514_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT119), .B(G141gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n851_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n851_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n858_), .A2(new_n717_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(G148gat), .Z(G1345gat));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n848_), .A2(new_n866_), .A3(new_n621_), .A4(new_n850_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT121), .B1(new_n858_), .B2(new_n622_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT61), .B(G155gat), .Z(new_n869_));
  AND3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1346gat));
  NAND4_X1  g671(.A1(new_n848_), .A2(new_n280_), .A3(new_n601_), .A4(new_n850_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G162gat), .B1(new_n858_), .B2(new_n668_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT122), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n873_), .A2(new_n874_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g678(.A1(new_n698_), .A2(new_n463_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n826_), .A2(new_n338_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n720_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  INV_X1    g683(.A(new_n882_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n357_), .A2(new_n358_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n218_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n887_), .B2(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(new_n717_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G176gat), .B1(new_n881_), .B2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT123), .B1(new_n833_), .B2(new_n338_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n857_), .A2(new_n893_), .A3(new_n464_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n220_), .B(new_n880_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n895_), .B2(new_n890_), .ZN(G1349gat));
  NOR2_X1   g695(.A1(new_n622_), .A2(new_n231_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n881_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n622_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n463_), .A3(new_n698_), .ZN(new_n900_));
  INV_X1    g699(.A(G183gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n881_), .A2(new_n361_), .A3(new_n601_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n881_), .A2(new_n606_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n233_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n647_), .A2(new_n454_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(KEYINPUT124), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n833_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n697_), .B1(KEYINPUT124), .B2(new_n906_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n720_), .A3(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n890_), .A3(new_n909_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n302_), .A2(KEYINPUT125), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n302_), .A2(KEYINPUT125), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT126), .Z(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OR3_X1    g715(.A1(new_n912_), .A2(new_n913_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1353gat));
  NAND2_X1  g718(.A1(new_n908_), .A2(new_n909_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT63), .B(G211gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n921_), .A2(new_n621_), .A3(new_n922_), .ZN(new_n923_));
  OAI22_X1  g722(.A1(new_n920_), .A2(new_n622_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n920_), .A2(new_n926_), .A3(new_n668_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n921_), .A2(new_n601_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1355gat));
endmodule


