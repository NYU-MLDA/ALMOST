//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT64), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G71gat), .B(G78gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n215_), .A2(new_n216_), .B1(new_n219_), .B2(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT8), .B1(new_n219_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n216_), .A3(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n231_), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n225_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n228_), .A2(new_n234_), .A3(new_n219_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  INV_X1    g035(.A(new_n218_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n227_), .A3(new_n238_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n234_), .A2(new_n219_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n226_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT66), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n226_), .B(new_n243_), .C1(new_n235_), .C2(new_n240_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n213_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n213_), .A3(new_n244_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n204_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n244_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n213_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT12), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G85gat), .B(G92gat), .ZN(new_n253_));
  OAI22_X1  g052(.A1(new_n221_), .A2(new_n253_), .B1(new_n214_), .B2(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n225_), .A2(new_n222_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n230_), .A2(new_n232_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n229_), .B2(new_n216_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n219_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n239_), .A2(new_n236_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n228_), .A2(new_n234_), .A3(new_n219_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n256_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT12), .B(new_n212_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n252_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n241_), .A2(KEYINPUT67), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n247_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n251_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n248_), .B1(new_n273_), .B2(new_n204_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n274_), .A2(new_n279_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n281_), .A2(KEYINPUT13), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT13), .B1(new_n281_), .B2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT73), .B(G1gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT74), .ZN(new_n293_));
  XOR2_X1   g092(.A(G1gat), .B(G8gat), .Z(new_n294_));
  OR2_X1    g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G29gat), .B(G36gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n297_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G229gat), .A2(G233gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n300_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n297_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n300_), .B(KEYINPUT15), .Z(new_n307_));
  NAND3_X1  g106(.A1(new_n295_), .A2(new_n296_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n302_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G113gat), .B(G141gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G169gat), .B(G197gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n304_), .B2(new_n310_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n287_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n316_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT79), .A3(new_n314_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n286_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT22), .B(G169gat), .ZN(new_n327_));
  INV_X1    g126(.A(G176gat), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT23), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT81), .B(G190gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n333_), .A2(G183gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n329_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(KEYINPUT26), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT25), .B(G183gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT80), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340_));
  INV_X1    g139(.A(G183gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(KEYINPUT25), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n336_), .A2(new_n337_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT24), .A3(new_n325_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n331_), .B(new_n346_), .C1(KEYINPUT24), .C2(new_n345_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n335_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n349_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G71gat), .B(G99gat), .ZN(new_n355_));
  INV_X1    g154(.A(G43gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G15gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n357_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT84), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n354_), .A2(new_n360_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT86), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT85), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G120gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT31), .Z(new_n372_));
  NOR2_X1   g171(.A1(new_n365_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n363_), .A2(KEYINPUT86), .A3(new_n364_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n363_), .A2(KEYINPUT86), .A3(new_n364_), .A4(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(KEYINPUT88), .A2(G141gat), .A3(G148gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(KEYINPUT3), .Z(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT2), .Z(new_n384_));
  OAI211_X1 g183(.A(new_n378_), .B(new_n380_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n378_), .A2(KEYINPUT1), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n378_), .B1(new_n379_), .B2(KEYINPUT1), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(KEYINPUT87), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(KEYINPUT87), .B2(new_n387_), .ZN(new_n389_));
  OR2_X1    g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n383_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT28), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G22gat), .B(G50gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  INV_X1    g198(.A(G228gat), .ZN(new_n400_));
  INV_X1    g199(.A(G233gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n393_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n405_), .A2(KEYINPUT21), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(KEYINPUT21), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G197gat), .B(G204gat), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n408_), .A3(KEYINPUT21), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n399_), .B(new_n402_), .C1(new_n404_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n403_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n392_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n402_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT92), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n393_), .A2(new_n394_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n411_), .B(KEYINPUT90), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n402_), .B(KEYINPUT89), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n418_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT93), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n422_), .A2(new_n419_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n428_), .B1(new_n413_), .B2(new_n417_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n425_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n398_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT94), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n432_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT95), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n423_), .A2(KEYINPUT95), .A3(new_n426_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n398_), .A4(new_n430_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n411_), .B(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n351_), .A3(new_n350_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(new_n326_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT99), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n344_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n445_), .B2(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n344_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT26), .B(G190gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n338_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n447_), .A2(new_n331_), .A3(new_n448_), .A4(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G183gat), .A2(G190gat), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n332_), .A2(KEYINPUT100), .A3(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT100), .B1(new_n332_), .B2(new_n452_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n329_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT101), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n411_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n456_), .B2(new_n411_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n442_), .B(KEYINPUT20), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT97), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT18), .ZN(new_n467_));
  XOR2_X1   g266(.A(G64gat), .B(G92gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n456_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n463_), .B1(new_n470_), .B2(new_n412_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n420_), .A2(new_n352_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT20), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n465_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n469_), .B1(new_n465_), .B2(new_n473_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G29gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT0), .ZN(new_n477_));
  INV_X1    g276(.A(G57gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G85gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n392_), .A2(new_n371_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n369_), .A2(new_n385_), .A3(new_n391_), .A4(new_n370_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G225gat), .A2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n483_), .A2(KEYINPUT4), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n489_), .A2(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(KEYINPUT4), .A3(new_n484_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT102), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT102), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n483_), .A2(new_n493_), .A3(KEYINPUT4), .A4(new_n484_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  AOI211_X1 g294(.A(new_n482_), .B(new_n488_), .C1(new_n490_), .C2(new_n495_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n474_), .A2(new_n475_), .A3(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n487_), .B1(new_n483_), .B2(KEYINPUT4), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT103), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n485_), .A2(new_n486_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(KEYINPUT33), .A3(new_n501_), .A4(new_n482_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT104), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n499_), .A2(KEYINPUT103), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT103), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n505_), .B(new_n498_), .C1(new_n492_), .C2(new_n494_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n501_), .B(new_n482_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT33), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n497_), .A2(new_n502_), .A3(new_n503_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n469_), .A2(KEYINPUT32), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n458_), .A2(new_n459_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n464_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(KEYINPUT20), .A3(new_n442_), .A4(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n470_), .A2(KEYINPUT105), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT105), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n456_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n411_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n472_), .A2(KEYINPUT20), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n463_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n511_), .B1(new_n514_), .B2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n465_), .A2(new_n473_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(new_n511_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n482_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n507_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n510_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n497_), .A2(new_n502_), .A3(new_n509_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT104), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n439_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n524_), .A2(new_n525_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n438_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n434_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT27), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n474_), .A2(KEYINPUT106), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n465_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT106), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n514_), .A2(new_n520_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n536_), .B(new_n539_), .C1(new_n469_), .C2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n535_), .B1(new_n541_), .B2(KEYINPUT27), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n534_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n377_), .B1(new_n530_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n377_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(new_n439_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n531_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n324_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n307_), .A2(new_n241_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n242_), .A2(new_n305_), .A3(new_n244_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n550_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n552_), .A2(new_n556_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT35), .B1(new_n557_), .B2(new_n560_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G190gat), .B(G218gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT71), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n570_), .A3(new_n567_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n566_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n213_), .B(new_n576_), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n297_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT75), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT76), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n584_), .B(KEYINPUT17), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n578_), .B2(KEYINPUT78), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(KEYINPUT78), .B2(new_n578_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n575_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n548_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n531_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT107), .Z(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n596_), .A2(KEYINPUT70), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(KEYINPUT70), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n599_));
  OAI22_X1  g398(.A1(new_n597_), .A2(new_n598_), .B1(new_n574_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n590_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n548_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n531_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n288_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT38), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n594_), .A2(new_n607_), .ZN(G1324gat));
  NAND3_X1  g407(.A1(new_n548_), .A2(new_n542_), .A3(new_n591_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(G8gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT108), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n609_), .A2(G8gat), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n613_), .B(new_n614_), .C1(new_n610_), .C2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n604_), .A2(new_n289_), .A3(new_n542_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n592_), .B2(new_n377_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT41), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT41), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n603_), .A2(G15gat), .A3(new_n377_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(new_n439_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G22gat), .B1(new_n592_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n626_), .A2(G22gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n603_), .B2(new_n629_), .ZN(G1327gat));
  INV_X1    g429(.A(new_n590_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n574_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n548_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n605_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n529_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n510_), .A2(new_n526_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n626_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n542_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n531_), .A3(new_n439_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n545_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  NOR4_X1   g440(.A1(new_n377_), .A2(new_n605_), .A3(new_n542_), .A4(new_n439_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n601_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT43), .B1(new_n643_), .B2(KEYINPUT110), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT110), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n600_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(KEYINPUT109), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n645_), .B(KEYINPUT43), .C1(new_n646_), .C2(KEYINPUT109), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n324_), .A2(new_n631_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n649_), .A4(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(G29gat), .A3(new_n605_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT109), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT110), .B1(new_n643_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n646_), .B2(new_n645_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n649_), .B(new_n650_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n635_), .B1(new_n652_), .B2(new_n659_), .ZN(G1328gat));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n651_), .A3(new_n542_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n633_), .A2(G36gat), .A3(new_n639_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT45), .Z(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(KEYINPUT46), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  NAND4_X1  g468(.A1(new_n659_), .A2(new_n651_), .A3(G43gat), .A4(new_n545_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n356_), .B1(new_n633_), .B2(new_n377_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT111), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g473(.A1(new_n659_), .A2(new_n439_), .A3(new_n651_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G50gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n626_), .A2(G50gat), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT112), .Z(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n633_), .B2(new_n678_), .ZN(G1331gat));
  INV_X1    g478(.A(new_n322_), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n680_), .B(new_n285_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n602_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n531_), .B1(new_n682_), .B2(KEYINPUT113), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(KEYINPUT113), .B2(new_n682_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n591_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n605_), .A2(KEYINPUT114), .A3(G57gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(KEYINPUT114), .B2(G57gat), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n684_), .A2(new_n478_), .B1(new_n686_), .B2(new_n688_), .ZN(G1332gat));
  OAI21_X1  g488(.A(G64gat), .B1(new_n685_), .B2(new_n639_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT48), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n639_), .A2(G64gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n682_), .B2(new_n692_), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n685_), .B2(new_n377_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n377_), .A2(G71gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n682_), .B2(new_n697_), .ZN(G1334gat));
  INV_X1    g497(.A(KEYINPUT50), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n686_), .A2(new_n439_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G78gat), .ZN(new_n701_));
  INV_X1    g500(.A(G78gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT50), .B(new_n702_), .C1(new_n686_), .C2(new_n439_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n439_), .A2(new_n702_), .ZN(new_n704_));
  OAI22_X1  g503(.A1(new_n701_), .A2(new_n703_), .B1(new_n682_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT116), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1335gat));
  NAND3_X1  g506(.A1(new_n286_), .A2(new_n322_), .A3(new_n590_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT117), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n648_), .A2(new_n649_), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n531_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n681_), .A2(new_n632_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n480_), .A3(new_n605_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1336gat));
  OAI21_X1  g514(.A(G92gat), .B1(new_n710_), .B2(new_n639_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n639_), .A2(G92gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n712_), .B2(new_n717_), .ZN(G1337gat));
  OAI21_X1  g517(.A(G99gat), .B1(new_n710_), .B2(new_n377_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n713_), .A2(new_n215_), .A3(new_n545_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n216_), .A3(new_n439_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n648_), .A2(new_n439_), .A3(new_n649_), .A4(new_n709_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(new_n725_), .A3(G106gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G106gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n723_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1339gat));
  NAND4_X1  g531(.A1(new_n600_), .A2(new_n322_), .A3(new_n285_), .A4(new_n631_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT54), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT122), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n273_), .B2(new_n204_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n247_), .B(new_n271_), .C1(new_n245_), .C2(KEYINPUT12), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(KEYINPUT55), .A3(new_n203_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT118), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n739_), .A2(new_n741_), .A3(new_n203_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n739_), .B2(new_n203_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n738_), .A2(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT119), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n739_), .A2(new_n203_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT118), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n739_), .A2(new_n741_), .A3(new_n203_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n251_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n272_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n737_), .A4(new_n204_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT55), .B1(new_n739_), .B2(new_n203_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(KEYINPUT119), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n279_), .B1(new_n746_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n736_), .B1(new_n757_), .B2(KEYINPUT56), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n750_), .A2(KEYINPUT119), .A3(new_n755_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT119), .B1(new_n750_), .B2(new_n755_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n278_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(KEYINPUT122), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n757_), .A2(KEYINPUT56), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n306_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n313_), .B(new_n767_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT120), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n769_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n319_), .A3(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n281_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n766_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n766_), .B1(new_n765_), .B2(new_n773_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n601_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n281_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n757_), .A2(KEYINPUT56), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n762_), .B(new_n279_), .C1(new_n746_), .C2(new_n756_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n281_), .A2(new_n282_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n772_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n575_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(KEYINPUT121), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n784_), .B2(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n784_), .A2(KEYINPUT57), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n777_), .A2(new_n787_), .A3(new_n789_), .A4(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n735_), .B1(new_n791_), .B2(new_n590_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n545_), .A2(new_n546_), .A3(new_n605_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT59), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT123), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n777_), .B(new_n795_), .C1(KEYINPUT57), .C2(new_n784_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n765_), .A2(new_n773_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT58), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n600_), .B1(new_n798_), .B2(new_n774_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n784_), .A2(KEYINPUT57), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT123), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n796_), .A2(new_n801_), .A3(new_n790_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n735_), .B1(new_n802_), .B2(new_n590_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n793_), .A2(KEYINPUT59), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n794_), .B(new_n680_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(G113gat), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n792_), .A2(new_n793_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n680_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT124), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n812_), .A3(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1340gat));
  OAI21_X1  g613(.A(new_n794_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G120gat), .B1(new_n815_), .B2(new_n285_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n817_));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n286_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n807_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(G1341gat));
  OAI21_X1  g621(.A(G127gat), .B1(new_n815_), .B2(new_n590_), .ZN(new_n823_));
  INV_X1    g622(.A(G127gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n807_), .A2(new_n824_), .A3(new_n631_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1342gat));
  OAI21_X1  g625(.A(G134gat), .B1(new_n815_), .B2(new_n600_), .ZN(new_n827_));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n807_), .A2(new_n828_), .A3(new_n575_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1343gat));
  INV_X1    g629(.A(new_n792_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n377_), .A2(new_n439_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(new_n531_), .A3(new_n542_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n322_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT125), .B(G141gat), .Z(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1344gat));
  INV_X1    g636(.A(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n286_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n631_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  OR3_X1    g642(.A1(new_n834_), .A2(G162gat), .A3(new_n574_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G162gat), .B1(new_n834_), .B2(new_n600_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1347gat));
  INV_X1    g645(.A(KEYINPUT126), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n377_), .A2(new_n639_), .A3(new_n605_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n626_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n790_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n798_), .A2(new_n774_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n800_), .B1(new_n852_), .B2(new_n601_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n853_), .B2(new_n795_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n631_), .B1(new_n854_), .B2(new_n801_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n680_), .B(new_n850_), .C1(new_n855_), .C2(new_n735_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n803_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n858_), .A2(new_n680_), .A3(new_n327_), .A4(new_n850_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT62), .B1(new_n856_), .B2(G169gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n847_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(G169gat), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT126), .A3(new_n857_), .A4(new_n859_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n866_), .ZN(G1348gat));
  NAND3_X1  g666(.A1(new_n848_), .A2(G176gat), .A3(new_n286_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n792_), .A2(new_n439_), .A3(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n803_), .A2(new_n849_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n286_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n871_), .B2(new_n328_), .ZN(G1349gat));
  NOR2_X1   g671(.A1(new_n590_), .A2(new_n338_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n831_), .A2(new_n626_), .A3(new_n631_), .A4(new_n848_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n870_), .A2(new_n873_), .B1(new_n874_), .B2(new_n341_), .ZN(G1350gat));
  NAND3_X1  g674(.A1(new_n870_), .A2(new_n449_), .A3(new_n575_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n803_), .A2(new_n600_), .A3(new_n849_), .ZN(new_n877_));
  INV_X1    g676(.A(G190gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1351gat));
  INV_X1    g678(.A(G197gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n832_), .A2(new_n639_), .A3(new_n605_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n831_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n882_), .B2(new_n322_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT127), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(KEYINPUT127), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n882_), .A2(new_n880_), .A3(new_n322_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(G1352gat));
  INV_X1    g686(.A(new_n882_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n286_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g689(.A1(new_n882_), .A2(new_n590_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n891_), .B2(new_n892_), .ZN(G1354gat));
  OR3_X1    g694(.A1(new_n882_), .A2(G218gat), .A3(new_n574_), .ZN(new_n896_));
  OAI21_X1  g695(.A(G218gat), .B1(new_n882_), .B2(new_n600_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1355gat));
endmodule


