//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT22), .B(G169gat), .Z(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT85), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT85), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n206_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n204_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n207_), .A2(new_n211_), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n219_), .C1(KEYINPUT24), .C2(new_n218_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n205_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT25), .B(G183gat), .Z(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(KEYINPUT83), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(new_n206_), .A3(KEYINPUT26), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT26), .B(G190gat), .Z(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(new_n224_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n220_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n214_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT86), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G211gat), .B(G218gat), .Z(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT94), .B(G197gat), .Z(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(G197gat), .B2(G204gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n232_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  MUX2_X1   g037(.A(G197gat), .B(new_n233_), .S(G204gat), .Z(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(KEYINPUT21), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT21), .A3(new_n232_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT20), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n215_), .A2(new_n213_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n204_), .B1(new_n246_), .B2(KEYINPUT98), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(KEYINPUT98), .B2(new_n246_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n202_), .A3(new_n218_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n222_), .A2(new_n226_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n212_), .A2(new_n251_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n245_), .A2(KEYINPUT96), .B1(new_n242_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(KEYINPUT96), .B2(new_n245_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G226gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT19), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT99), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n231_), .A2(new_n243_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n255_), .B2(new_n242_), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n263_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT18), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n262_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n259_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n263_), .A2(new_n277_), .A3(new_n264_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n257_), .B2(new_n277_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n275_), .B1(new_n279_), .B2(new_n271_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G127gat), .B(G134gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT89), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT90), .ZN(new_n285_));
  XOR2_X1   g084(.A(G113gat), .B(G120gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(G141gat), .ZN(new_n289_));
  INV_X1    g088(.A(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(KEYINPUT92), .A3(KEYINPUT1), .ZN(new_n293_));
  OR2_X1    g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n293_), .B(new_n294_), .C1(KEYINPUT1), .C2(new_n292_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT92), .B1(new_n292_), .B2(KEYINPUT1), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n288_), .B(new_n291_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n288_), .B(KEYINPUT2), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n291_), .A2(KEYINPUT3), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n291_), .A2(KEYINPUT3), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT93), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n294_), .A2(new_n292_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n297_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n287_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n287_), .A2(new_n304_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n305_), .A2(KEYINPUT4), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n287_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n307_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n305_), .A2(new_n306_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(new_n311_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G29gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT0), .ZN(new_n316_));
  INV_X1    g115(.A(G57gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G85gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n314_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n243_), .B1(new_n304_), .B2(KEYINPUT29), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(KEYINPUT95), .B2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(KEYINPUT95), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n304_), .A2(KEYINPUT29), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT28), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n334_), .B(new_n336_), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n231_), .B(KEYINPUT30), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G15gat), .B(G43gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n339_), .B(KEYINPUT87), .Z(new_n340_));
  XOR2_X1   g139(.A(G71gat), .B(G99gat), .Z(new_n341_));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n340_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n338_), .B(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT91), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n287_), .B(KEYINPUT31), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n350_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n337_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n334_), .B(new_n336_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n353_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n282_), .B(new_n325_), .C1(new_n356_), .C2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n323_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT33), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(KEYINPUT33), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n309_), .A2(new_n311_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n313_), .B(KEYINPUT101), .Z(new_n365_));
  OAI221_X1 g164(.A(new_n320_), .B1(new_n307_), .B2(new_n364_), .C1(new_n365_), .C2(new_n311_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n266_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n279_), .A2(new_n368_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n324_), .A2(new_n370_), .ZN(new_n371_));
  OAI22_X1  g170(.A1(new_n367_), .A2(new_n274_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n360_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G230gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(G106gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT64), .B1(new_n382_), .B2(new_n377_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n376_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G85gat), .A2(G92gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G85gat), .A2(G92gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n387_), .B2(KEYINPUT9), .ZN(new_n388_));
  INV_X1    g187(.A(G92gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT65), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G92gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n319_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n388_), .B1(new_n393_), .B2(KEYINPUT9), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G99gat), .A2(G106gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT6), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n384_), .A2(new_n394_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n384_), .A2(new_n394_), .A3(KEYINPUT66), .A4(new_n400_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n405_));
  INV_X1    g204(.A(G99gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n376_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT67), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT7), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT7), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT67), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n408_), .A2(new_n406_), .A3(new_n376_), .A4(KEYINPUT7), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n399_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n385_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT8), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n386_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n405_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  OAI22_X1  g217(.A1(new_n410_), .A2(KEYINPUT67), .B1(G99gat), .B2(G106gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n408_), .A2(KEYINPUT7), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n413_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n400_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n417_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT68), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT69), .B1(new_n397_), .B2(new_n398_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n397_), .A2(KEYINPUT69), .A3(new_n398_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n421_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n415_), .A2(new_n386_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n416_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n403_), .B(new_n404_), .C1(new_n425_), .C2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT70), .B(G71gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G78gat), .ZN(new_n436_));
  INV_X1    g235(.A(G78gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G57gat), .B(G64gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT11), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n439_), .A2(KEYINPUT11), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n436_), .B(new_n438_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n438_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n434_), .A2(new_n437_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n440_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n375_), .B1(new_n433_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT69), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(new_n426_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n430_), .B1(new_n456_), .B2(new_n421_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n418_), .B(new_n424_), .C1(new_n457_), .C2(new_n416_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(new_n404_), .A3(new_n403_), .A4(new_n447_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT72), .A3(new_n375_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n433_), .B2(new_n448_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n433_), .A2(new_n461_), .A3(new_n448_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n451_), .B(new_n460_), .C1(new_n462_), .C2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n459_), .A2(KEYINPUT71), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n403_), .A2(new_n404_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT71), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n458_), .A4(new_n447_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n433_), .A2(new_n448_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n375_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G120gat), .B(G148gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT5), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G176gat), .B(G204gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n465_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT74), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n465_), .A2(new_n473_), .A3(new_n480_), .A4(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n459_), .A2(KEYINPUT72), .A3(new_n375_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT72), .B1(new_n459_), .B2(new_n375_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n462_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n463_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n485_), .A2(new_n487_), .B1(new_n472_), .B2(new_n471_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n477_), .B(KEYINPUT73), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n482_), .A2(KEYINPUT13), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT13), .B1(new_n482_), .B2(new_n491_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G113gat), .B(G141gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT82), .ZN(new_n497_));
  XOR2_X1   g296(.A(G169gat), .B(G197gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G22gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G15gat), .ZN(new_n501_));
  INV_X1    g300(.A(G15gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G22gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G1gat), .A2(G8gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n505_), .A2(KEYINPUT14), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT78), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT78), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(KEYINPUT14), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G1gat), .ZN(new_n512_));
  INV_X1    g311(.A(G8gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n505_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT79), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(new_n517_), .A3(new_n505_), .ZN(new_n518_));
  AND4_X1   g317(.A1(new_n507_), .A2(new_n511_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n507_), .A2(new_n511_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n520_));
  INV_X1    g319(.A(G36gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(G29gat), .ZN(new_n522_));
  INV_X1    g321(.A(G29gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G36gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G43gat), .ZN(new_n526_));
  INV_X1    g325(.A(G50gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G43gat), .A2(G50gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n528_), .A2(new_n522_), .A3(new_n524_), .A4(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n519_), .A2(new_n520_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n507_), .A2(new_n511_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n516_), .A2(new_n518_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n507_), .A2(new_n511_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n533_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n535_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n534_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n533_), .A2(KEYINPUT15), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT15), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n531_), .A2(new_n532_), .A3(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n538_), .A2(new_n545_), .A3(new_n539_), .A4(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n499_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n542_), .A2(new_n549_), .A3(new_n499_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n495_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n374_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT80), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n447_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n538_), .A2(new_n539_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT16), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n560_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n565_), .B(KEYINPUT17), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n545_), .A2(new_n547_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n433_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  OAI221_X1 g374(.A(new_n573_), .B1(KEYINPUT35), .B2(new_n575_), .C1(new_n433_), .C2(new_n533_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT75), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n579_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT36), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT77), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n576_), .B(new_n578_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(KEYINPUT77), .A3(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n580_), .A2(new_n581_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n588_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n571_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n555_), .A2(new_n324_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G1gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n586_), .A2(KEYINPUT76), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n600_), .A3(new_n585_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n601_), .A3(new_n593_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n588_), .A2(new_n590_), .A3(new_n593_), .A4(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n571_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n555_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n512_), .A3(new_n324_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n598_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n612_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT102), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(G1324gat));
  INV_X1    g420(.A(new_n282_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n610_), .A2(new_n513_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n555_), .A2(new_n596_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G8gat), .B1(new_n624_), .B2(new_n282_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n624_), .B2(new_n354_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT41), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n610_), .A2(new_n502_), .A3(new_n353_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(G1326gat));
  XOR2_X1   g433(.A(new_n357_), .B(KEYINPUT104), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G22gat), .B1(new_n624_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT42), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n610_), .A2(new_n500_), .A3(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n607_), .A2(new_n594_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n555_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n324_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n554_), .A2(new_n571_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n606_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n374_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT43), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n374_), .A2(new_n648_), .A3(new_n645_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n644_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT44), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n652_), .A2(new_n523_), .A3(new_n325_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n650_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(KEYINPUT105), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n650_), .B2(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n643_), .B1(new_n653_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n651_), .A2(new_n622_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n521_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n642_), .A2(new_n521_), .A3(new_n622_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n661_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n658_), .B2(new_n656_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT46), .B(new_n666_), .C1(new_n669_), .C2(new_n521_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1329gat));
  AOI21_X1  g470(.A(G43gat), .B1(new_n642_), .B2(new_n353_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n526_), .B(new_n354_), .C1(new_n650_), .C2(KEYINPUT44), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n659_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1330gat));
  AOI21_X1  g475(.A(G50gat), .B1(new_n642_), .B2(new_n635_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n652_), .A2(new_n527_), .A3(new_n357_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n659_), .ZN(G1331gat));
  INV_X1    g478(.A(new_n553_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n494_), .A2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n374_), .A2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(new_n609_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n596_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n325_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1332gat));
  OAI21_X1  g486(.A(G64gat), .B1(new_n685_), .B2(new_n282_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT48), .ZN(new_n689_));
  INV_X1    g488(.A(G64gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n690_), .A3(new_n622_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1333gat));
  OAI21_X1  g491(.A(G71gat), .B1(new_n685_), .B2(new_n354_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT49), .ZN(new_n694_));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n683_), .A2(new_n695_), .A3(new_n353_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1334gat));
  OAI21_X1  g496(.A(G78gat), .B1(new_n685_), .B2(new_n636_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT50), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n683_), .A2(new_n437_), .A3(new_n635_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1335gat));
  NAND2_X1  g500(.A1(new_n682_), .A2(new_n641_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n319_), .B1(new_n702_), .B2(new_n325_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT106), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n681_), .A2(new_n571_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n325_), .A2(new_n319_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(new_n389_), .B1(new_n702_), .B2(new_n282_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT107), .Z(new_n710_));
  AOI21_X1  g509(.A(new_n282_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n706_), .B2(new_n711_), .ZN(G1337gat));
  OAI21_X1  g511(.A(new_n353_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n702_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n706_), .A2(new_n353_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G99gat), .ZN(new_n716_));
  AND4_X1   g515(.A1(KEYINPUT108), .A2(new_n716_), .A3(KEYINPUT109), .A4(KEYINPUT51), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT51), .B1(new_n716_), .B2(KEYINPUT109), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(KEYINPUT108), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(G1338gat));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n706_), .A2(new_n337_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G106gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT52), .B(new_n376_), .C1(new_n706_), .C2(new_n337_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n337_), .A2(new_n376_), .ZN(new_n725_));
  OAI22_X1  g524(.A1(new_n723_), .A2(new_n724_), .B1(new_n702_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g526(.A(KEYINPUT120), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n608_), .A2(new_n495_), .A3(new_n680_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n544_), .A2(new_n548_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n544_), .A2(new_n548_), .A3(KEYINPUT114), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n541_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n541_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n499_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n732_), .B(new_n550_), .C1(new_n737_), .C2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n544_), .A2(new_n548_), .A3(KEYINPUT114), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT114), .B1(new_n544_), .B2(new_n548_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n543_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n738_), .A2(new_n739_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n732_), .B1(new_n747_), .B2(new_n550_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n742_), .A2(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT117), .B(new_n749_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n751_));
  INV_X1    g550(.A(new_n749_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n482_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n750_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n451_), .A2(new_n460_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n464_), .A2(new_n462_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT112), .B(new_n755_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n466_), .A2(new_n469_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n472_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n465_), .B2(KEYINPUT112), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n490_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT56), .B(new_n490_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT58), .B1(new_n754_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT118), .B1(new_n768_), .B2(new_n606_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n480_), .B1(new_n488_), .B2(new_n477_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n481_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n752_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT117), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n482_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n766_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT112), .B1(new_n756_), .B2(new_n757_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT55), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n780_), .B2(new_n490_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n770_), .B1(new_n776_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n645_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n754_), .A2(KEYINPUT58), .A3(new_n767_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n769_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n482_), .B2(new_n680_), .ZN(new_n790_));
  AOI211_X1 g589(.A(KEYINPUT111), .B(new_n553_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n765_), .A2(new_n793_), .A3(new_n766_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n780_), .A2(KEYINPUT113), .A3(KEYINPUT56), .A4(new_n490_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n482_), .A2(new_n491_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n752_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n594_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n594_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n788_), .A2(new_n802_), .A3(KEYINPUT119), .A4(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n571_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n774_), .B(new_n775_), .C1(new_n777_), .C2(new_n781_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n606_), .B1(new_n806_), .B2(new_n770_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n786_), .B1(new_n807_), .B2(new_n784_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n808_), .A2(new_n769_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT119), .B1(new_n809_), .B2(new_n803_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n728_), .B(new_n731_), .C1(new_n805_), .C2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n788_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n571_), .A3(new_n804_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n728_), .B1(new_n816_), .B2(new_n731_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n812_), .A2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n622_), .A2(new_n325_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n359_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n680_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n809_), .A2(KEYINPUT121), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n803_), .B1(new_n809_), .B2(KEYINPUT121), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n571_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n731_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n820_), .A2(KEYINPUT59), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n822_), .A2(KEYINPUT59), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n680_), .A2(new_n831_), .A3(G113gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n831_), .B2(G113gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n824_), .B1(new_n830_), .B2(new_n833_), .ZN(G1340gat));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n495_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n823_), .A2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n830_), .A2(new_n495_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n836_), .ZN(G1341gat));
  AND2_X1   g640(.A1(new_n830_), .A2(new_n607_), .ZN(new_n842_));
  INV_X1    g641(.A(G127gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n607_), .A2(new_n843_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n842_), .A2(new_n843_), .B1(new_n822_), .B2(new_n844_), .ZN(G1342gat));
  AOI21_X1  g644(.A(G134gat), .B1(new_n823_), .B2(new_n595_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT123), .B(G134gat), .Z(new_n847_));
  NOR2_X1   g646(.A1(new_n606_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n830_), .B2(new_n848_), .ZN(G1343gat));
  NAND3_X1  g648(.A1(new_n818_), .A2(new_n356_), .A3(new_n819_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n553_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(new_n289_), .ZN(G1344gat));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n494_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n290_), .ZN(G1345gat));
  NOR2_X1   g653(.A1(new_n850_), .A2(new_n571_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT61), .B(G155gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n850_), .B2(new_n606_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n594_), .A2(G162gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n850_), .B2(new_n859_), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n282_), .A2(new_n324_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n353_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n635_), .B(new_n862_), .C1(new_n827_), .C2(new_n731_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n680_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n203_), .B2(new_n864_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT62), .B1(new_n864_), .B2(G169gat), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1348gat));
  AOI21_X1  g667(.A(G176gat), .B1(new_n863_), .B2(new_n495_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n818_), .A2(new_n357_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT124), .Z(new_n871_));
  NOR3_X1   g670(.A1(new_n862_), .A2(new_n217_), .A3(new_n494_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  NAND4_X1  g672(.A1(new_n871_), .A2(new_n607_), .A3(new_n353_), .A4(new_n861_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n607_), .A2(new_n222_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n205_), .B1(new_n863_), .B2(new_n876_), .ZN(G1350gat));
  INV_X1    g676(.A(new_n226_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n863_), .A2(new_n595_), .A3(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n863_), .A2(new_n645_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n206_), .ZN(G1351gat));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n818_), .A2(new_n882_), .A3(new_n356_), .A4(new_n861_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n731_), .B1(new_n805_), .B2(new_n810_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT120), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n885_), .A2(new_n356_), .A3(new_n811_), .A4(new_n861_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n680_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n495_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g691(.A(new_n571_), .B1(new_n883_), .B2(new_n887_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n607_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT126), .B1(new_n900_), .B2(new_n894_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n893_), .A2(new_n902_), .A3(new_n895_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n897_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT127), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n897_), .B(new_n906_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1354gat));
  INV_X1    g707(.A(G218gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n888_), .A2(new_n909_), .A3(new_n595_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n606_), .B1(new_n883_), .B2(new_n887_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n909_), .ZN(G1355gat));
endmodule


