//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT64), .ZN(new_n203_));
  OAI211_X1 g002(.A(G85gat), .B(G92gat), .C1(KEYINPUT65), .C2(KEYINPUT9), .ZN(new_n204_));
  OAI211_X1 g003(.A(KEYINPUT65), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(G106gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n208_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n224_), .A2(KEYINPUT67), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT67), .B1(new_n224_), .B2(new_n225_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n213_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n217_), .B(new_n223_), .C1(new_n228_), .C2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n233_), .B(new_n213_), .C1(new_n227_), .C2(new_n226_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n217_), .B1(new_n237_), .B2(new_n223_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n216_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n223_), .B1(new_n228_), .B2(new_n234_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n217_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n235_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT69), .A3(new_n216_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n241_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n248_), .B1(new_n241_), .B2(new_n253_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n203_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n248_), .B(KEYINPUT70), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n256_), .B2(KEYINPUT12), .ZN(new_n260_));
  INV_X1    g059(.A(new_n203_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n257_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT5), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n257_), .B(new_n269_), .C1(new_n260_), .C2(new_n262_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n272_));
  NAND2_X1  g071(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n271_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G36gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G29gat), .ZN(new_n280_));
  INV_X1    g079(.A(G29gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G36gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G50gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G43gat), .ZN(new_n285_));
  INV_X1    g084(.A(G43gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G50gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G29gat), .B(G36gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G43gat), .B(G50gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n241_), .A2(new_n294_), .A3(new_n253_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n283_), .A2(new_n288_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n291_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT15), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT15), .B1(new_n296_), .B2(new_n297_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT35), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G232gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT34), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n239_), .A2(new_n301_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n295_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(new_n302_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G190gat), .B(G218gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G134gat), .B(G162gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(KEYINPUT36), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n308_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n313_), .B(KEYINPUT36), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT37), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n315_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n318_), .B1(new_n322_), .B2(new_n309_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT37), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n316_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT14), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(G1gat), .B2(G8gat), .ZN(new_n328_));
  INV_X1    g127(.A(G15gat), .ZN(new_n329_));
  INV_X1    g128(.A(G22gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G15gat), .A2(G22gat), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n328_), .A2(KEYINPUT72), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n334_));
  AND2_X1   g133(.A1(G1gat), .A2(G8gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n327_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G1gat), .A2(G8gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT73), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(G1gat), .A2(G8gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G1gat), .A2(G8gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n333_), .A2(new_n336_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(new_n332_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n336_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n338_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G231gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(new_n258_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G127gat), .B(G155gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(G183gat), .B(G211gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n354_), .A3(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(KEYINPUT17), .Z(new_n361_));
  INV_X1    g160(.A(new_n248_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n351_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n351_), .A2(new_n362_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n326_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT76), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT23), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(G169gat), .ZN(new_n375_));
  INV_X1    g174(.A(G176gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n373_), .B(new_n374_), .C1(new_n377_), .C2(KEYINPUT24), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT24), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT90), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n383_), .A3(KEYINPUT24), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n377_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  INV_X1    g186(.A(G183gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT25), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G183gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n385_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n386_), .B1(new_n385_), .B2(new_n392_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n379_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n373_), .B(new_n374_), .C1(G183gat), .C2(G190gat), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n396_), .A2(new_n380_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT22), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G169gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n375_), .A2(KEYINPUT22), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n397_), .B1(G176gat), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G197gat), .A2(G204gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT21), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(KEYINPUT21), .A3(new_n405_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n403_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT19), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT22), .B1(new_n375_), .B2(KEYINPUT84), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n376_), .C1(KEYINPUT84), .C2(new_n399_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n421_), .A2(new_n396_), .A3(new_n380_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n377_), .A2(KEYINPUT24), .A3(new_n380_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n388_), .B2(KEYINPUT25), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n390_), .A2(KEYINPUT82), .A3(G183gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT26), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT26), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G190gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n431_), .A3(new_n389_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n423_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n378_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT83), .B(new_n423_), .C1(new_n427_), .C2(new_n432_), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n419_), .B(new_n422_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(new_n379_), .A3(new_n436_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n422_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT85), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n413_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n418_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n440_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n419_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n413_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n439_), .A2(KEYINPUT85), .A3(new_n440_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n403_), .B2(new_n413_), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT92), .B(new_n447_), .C1(new_n395_), .C2(new_n402_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n449_), .B(KEYINPUT20), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n417_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT93), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n456_), .A3(new_n417_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n444_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT18), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G64gat), .B(G92gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  NOR2_X1   g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n453_), .A2(new_n456_), .A3(new_n417_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n456_), .B1(new_n453_), .B2(new_n417_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n462_), .B(new_n443_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n370_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n470_), .A2(G228gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(G228gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G78gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G22gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n479_));
  INV_X1    g278(.A(G141gat), .ZN(new_n480_));
  INV_X1    g279(.A(G148gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G141gat), .A2(G148gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G155gat), .B(G162gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(KEYINPUT1), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(KEYINPUT1), .B2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n480_), .A2(new_n481_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n483_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n499_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT28), .B1(new_n499_), .B2(KEYINPUT29), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n447_), .B1(new_n499_), .B2(KEYINPUT29), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n478_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n506_), .A3(new_n478_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n511_));
  NAND3_X1  g310(.A1(new_n446_), .A2(KEYINPUT30), .A3(new_n448_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(new_n329_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G71gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(G99gat), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n512_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n511_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G127gat), .B(G134gat), .Z(new_n523_));
  XOR2_X1   g322(.A(G113gat), .B(G120gat), .Z(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT86), .B(G43gat), .Z(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  NOR3_X1   g326(.A1(new_n437_), .A2(new_n441_), .A3(new_n513_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT30), .B1(new_n446_), .B2(new_n448_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n518_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n511_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n512_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n522_), .A2(new_n527_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n527_), .B1(new_n522_), .B2(new_n533_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n510_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n527_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n520_), .A2(new_n521_), .A3(new_n511_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n504_), .A2(new_n506_), .A3(new_n478_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n507_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n522_), .A2(new_n533_), .A3(new_n527_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n403_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n395_), .A2(KEYINPUT96), .A3(new_n402_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n447_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n442_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT97), .B1(new_n549_), .B2(KEYINPUT20), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n417_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n453_), .A2(new_n417_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n462_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT27), .A3(new_n466_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n499_), .A2(new_n525_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n525_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n492_), .A2(new_n561_), .A3(new_n498_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(KEYINPUT4), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT4), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n499_), .A2(new_n564_), .A3(new_n525_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G225gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT94), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G29gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G85gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT0), .B(G57gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT98), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n580_), .A3(new_n575_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n468_), .A2(new_n545_), .A3(new_n559_), .A4(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n443_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n557_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n560_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n586_), .A2(new_n573_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT95), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n563_), .A2(new_n566_), .A3(new_n565_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(KEYINPUT95), .B2(new_n587_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n575_), .A2(KEYINPUT33), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n568_), .A2(new_n592_), .A3(new_n569_), .A4(new_n574_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n588_), .A2(new_n590_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n466_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n579_), .A2(new_n575_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n443_), .B(new_n597_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n549_), .A2(KEYINPUT20), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n442_), .A3(new_n550_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n554_), .B1(new_n602_), .B2(new_n417_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n596_), .B(new_n598_), .C1(new_n603_), .C2(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n534_), .A2(new_n535_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n510_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n583_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n610_));
  XOR2_X1   g409(.A(G113gat), .B(G141gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT79), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n343_), .A2(new_n348_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(new_n294_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT77), .B1(new_n301_), .B2(new_n349_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT15), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n621_), .A2(new_n343_), .A3(new_n348_), .A4(new_n298_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT77), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n618_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n349_), .A2(new_n293_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n617_), .A2(new_n294_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n616_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT78), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n614_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n625_), .A2(KEYINPUT78), .A3(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT80), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n615_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n622_), .A2(new_n623_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n301_), .A2(new_n349_), .A3(KEYINPUT77), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n615_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n631_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n614_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n640_), .A2(new_n633_), .A3(KEYINPUT80), .A4(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n625_), .A2(new_n629_), .A3(new_n613_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT81), .B1(new_n634_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n640_), .A2(new_n633_), .A3(new_n641_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT80), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT81), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n643_), .A4(new_n642_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n609_), .A2(new_n610_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n585_), .A2(new_n466_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n370_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n653_), .A2(new_n370_), .B1(new_n654_), .B2(new_n558_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n582_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n536_), .B2(new_n544_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n655_), .A2(new_n657_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n651_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT99), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n278_), .B(new_n369_), .C1(new_n652_), .C2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT100), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(KEYINPUT100), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n582_), .A2(G1gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n664_), .A2(KEYINPUT38), .A3(new_n665_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n317_), .A2(new_n320_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n658_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT101), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n277_), .A2(new_n651_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(new_n366_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n582_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n668_), .A2(new_n669_), .A3(new_n677_), .ZN(G1324gat));
  NOR2_X1   g477(.A1(new_n655_), .A2(G8gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n662_), .A2(new_n663_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n655_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n672_), .A2(new_n681_), .A3(new_n674_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G8gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G8gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1325gat));
  NAND3_X1  g487(.A1(new_n661_), .A2(new_n329_), .A3(new_n606_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n672_), .A2(new_n606_), .A3(new_n674_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n690_), .B2(G15gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT102), .Z(G1326gat));
  XNOR2_X1  g493(.A(new_n510_), .B(KEYINPUT103), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n661_), .A2(new_n330_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n695_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G22gat), .B1(new_n676_), .B2(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(KEYINPUT42), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(KEYINPUT42), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(G1327gat));
  NAND3_X1  g500(.A1(new_n277_), .A2(new_n366_), .A3(new_n670_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n660_), .B2(new_n652_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G29gat), .B1(new_n703_), .B2(new_n656_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n658_), .B2(new_n326_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  INV_X1    g505(.A(new_n326_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n609_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n277_), .A2(new_n651_), .A3(new_n366_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT44), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n713_), .B(new_n710_), .C1(new_n705_), .C2(new_n708_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n582_), .A2(new_n281_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n704_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  AOI21_X1  g516(.A(new_n706_), .B1(new_n609_), .B2(new_n707_), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT43), .B(new_n326_), .C1(new_n583_), .C2(new_n608_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n711_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n713_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n709_), .A2(KEYINPUT44), .A3(new_n711_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n681_), .A3(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n655_), .A2(G36gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n703_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT45), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT104), .B1(new_n723_), .B2(G36gat), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT105), .B(KEYINPUT46), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n712_), .A2(new_n714_), .A3(new_n655_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n279_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n724_), .A3(new_n727_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT46), .B1(new_n735_), .B2(KEYINPUT105), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n731_), .A2(new_n736_), .ZN(G1329gat));
  AOI21_X1  g536(.A(G43gat), .B1(new_n703_), .B2(new_n606_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n606_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n286_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n715_), .B2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g541(.A1(new_n703_), .A2(new_n284_), .A3(new_n695_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n712_), .A2(new_n714_), .A3(new_n542_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT106), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n284_), .B1(new_n744_), .B2(KEYINPUT106), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n748_), .B2(new_n749_), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n277_), .A2(new_n651_), .A3(new_n366_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n672_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n582_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n369_), .A2(new_n277_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n658_), .A2(new_n651_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n656_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n757_), .B2(new_n759_), .ZN(G1332gat));
  OR3_X1    g559(.A1(new_n757_), .A2(G64gat), .A3(new_n655_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G64gat), .B1(new_n753_), .B2(new_n655_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT48), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT48), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1333gat));
  OR3_X1    g564(.A1(new_n757_), .A2(G71gat), .A3(new_n739_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G71gat), .B1(new_n753_), .B2(new_n739_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT49), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT49), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(G1334gat));
  OR3_X1    g569(.A1(new_n757_), .A2(G78gat), .A3(new_n697_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G78gat), .B1(new_n753_), .B2(new_n697_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT50), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT50), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(G1335gat));
  INV_X1    g574(.A(new_n670_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n277_), .A2(new_n367_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n756_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n218_), .A3(new_n656_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n277_), .A2(new_n651_), .A3(new_n367_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n709_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n656_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n783_), .B2(new_n218_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT108), .ZN(G1336gat));
  NAND3_X1  g584(.A1(new_n779_), .A2(new_n219_), .A3(new_n681_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n782_), .A2(new_n681_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n219_), .ZN(G1337gat));
  NOR3_X1   g587(.A1(new_n778_), .A2(new_n739_), .A3(new_n214_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n606_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G99gat), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT109), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n792_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT110), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n779_), .A2(new_n475_), .A3(new_n510_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n709_), .A2(new_n510_), .A3(new_n781_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT111), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n475_), .B1(new_n799_), .B2(KEYINPUT111), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n798_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT53), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n798_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1339gat));
  AOI22_X1  g608(.A1(new_n275_), .A2(new_n276_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n651_), .A2(new_n366_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n270_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n616_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n613_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n627_), .B(new_n616_), .C1(new_n619_), .C2(new_n624_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n817_), .B2(new_n613_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(KEYINPUT113), .A3(new_n643_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT113), .B1(new_n822_), .B2(new_n643_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n816_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n254_), .A2(new_n261_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT69), .B1(new_n252_), .B2(new_n216_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n208_), .A2(new_n215_), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n240_), .B(new_n831_), .C1(new_n251_), .C2(new_n235_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n362_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT12), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n829_), .A2(new_n835_), .A3(KEYINPUT55), .A4(new_n259_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n254_), .B(new_n259_), .C1(new_n256_), .C2(KEYINPUT12), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n203_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n828_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n839_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n839_), .B2(new_n267_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n826_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n326_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n826_), .B(KEYINPUT58), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n267_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT56), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n839_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n852_), .A2(KEYINPUT114), .A3(KEYINPUT58), .A4(new_n826_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n844_), .A2(new_n847_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n268_), .A2(new_n270_), .B1(new_n825_), .B2(new_n823_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n816_), .B1(new_n645_), .B2(new_n650_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n852_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n858_), .B2(new_n670_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n856_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n776_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n854_), .A2(new_n859_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n815_), .B1(new_n864_), .B2(new_n366_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n655_), .A2(new_n656_), .A3(new_n542_), .A4(new_n606_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n651_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n868_), .A2(KEYINPUT115), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(KEYINPUT115), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n866_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n866_), .A2(KEYINPUT116), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n866_), .A2(KEYINPUT116), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n862_), .B2(new_n776_), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n855_), .B(new_n670_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n367_), .B1(new_n878_), .B2(new_n854_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n879_), .B2(new_n815_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n871_), .A2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n651_), .A2(G113gat), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n869_), .A2(new_n870_), .B1(new_n881_), .B2(new_n882_), .ZN(G1340gat));
  NAND3_X1  g682(.A1(new_n871_), .A2(new_n880_), .A3(new_n278_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT117), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n871_), .A2(new_n880_), .A3(new_n886_), .A4(new_n278_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(G120gat), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n277_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n867_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n889_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT118), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n888_), .A2(new_n894_), .A3(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1341gat));
  AOI21_X1  g695(.A(G127gat), .B1(new_n867_), .B2(new_n367_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n366_), .A2(KEYINPUT119), .ZN(new_n898_));
  MUX2_X1   g697(.A(KEYINPUT119), .B(new_n898_), .S(G127gat), .Z(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n881_), .B2(new_n899_), .ZN(G1342gat));
  INV_X1    g699(.A(G134gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n867_), .A2(new_n901_), .A3(new_n670_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n881_), .A2(new_n707_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n901_), .ZN(G1343gat));
  NOR2_X1   g703(.A1(new_n865_), .A2(new_n536_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n681_), .A2(new_n582_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n659_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT120), .B(G141gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1344gat));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n277_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n481_), .ZN(G1345gat));
  OR3_X1    g711(.A1(new_n907_), .A2(KEYINPUT121), .A3(new_n366_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT121), .B1(new_n907_), .B2(new_n366_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n915_), .B(new_n917_), .ZN(G1346gat));
  OR3_X1    g717(.A1(new_n907_), .A2(G162gat), .A3(new_n776_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G162gat), .B1(new_n907_), .B2(new_n326_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1347gat));
  INV_X1    g720(.A(new_n865_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n655_), .A2(new_n656_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n606_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT122), .B1(new_n924_), .B2(new_n659_), .ZN(new_n925_));
  OR3_X1    g724(.A1(new_n924_), .A2(KEYINPUT122), .A3(new_n659_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n922_), .A2(new_n697_), .A3(new_n925_), .A4(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(G169gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT123), .B1(new_n928_), .B2(KEYINPUT62), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(KEYINPUT62), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n927_), .A2(new_n931_), .A3(new_n932_), .A4(G169gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n929_), .A2(new_n930_), .A3(new_n933_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n865_), .A2(new_n695_), .A3(new_n924_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n659_), .A2(new_n401_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT124), .Z(new_n938_));
  OAI21_X1  g737(.A(new_n934_), .B1(new_n936_), .B2(new_n938_), .ZN(G1348gat));
  NAND2_X1  g738(.A1(new_n922_), .A2(new_n542_), .ZN(new_n940_));
  NOR4_X1   g739(.A1(new_n940_), .A2(new_n376_), .A3(new_n277_), .A4(new_n924_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G176gat), .B1(new_n935_), .B2(new_n278_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n942_), .A2(KEYINPUT125), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(KEYINPUT125), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n943_), .B2(new_n944_), .ZN(G1349gat));
  OR3_X1    g744(.A1(new_n940_), .A2(new_n366_), .A3(new_n924_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n366_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n946_), .A2(new_n388_), .B1(new_n935_), .B2(new_n947_), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n936_), .B2(new_n326_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n935_), .A2(new_n387_), .A3(new_n670_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1351gat));
  XOR2_X1   g750(.A(KEYINPUT126), .B(G197gat), .Z(new_n952_));
  NOR2_X1   g751(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n905_), .A2(new_n923_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n659_), .ZN(new_n955_));
  MUX2_X1   g754(.A(new_n952_), .B(new_n953_), .S(new_n955_), .Z(G1352gat));
  INV_X1    g755(.A(new_n954_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n278_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n367_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  AND2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n960_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n963_), .B1(new_n960_), .B2(new_n961_), .ZN(G1354gat));
  AOI21_X1  g763(.A(G218gat), .B1(new_n957_), .B2(new_n670_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n707_), .A2(G218gat), .ZN(new_n966_));
  XOR2_X1   g765(.A(new_n966_), .B(KEYINPUT127), .Z(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n957_), .B2(new_n967_), .ZN(G1355gat));
endmodule


