//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_;
  INV_X1    g000(.A(G57gat), .ZN(new_n202_));
  INV_X1    g001(.A(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n210_), .A3(new_n205_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G127gat), .B(G155gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G183gat), .B(G211gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT73), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222_));
  INV_X1    g021(.A(G1gat), .ZN(new_n223_));
  INV_X1    g022(.A(G8gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G1gat), .B(G8gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G231gat), .ZN(new_n231_));
  INV_X1    g030(.A(G233gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(KEYINPUT73), .B(new_n228_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n230_), .B2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n214_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n238_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n214_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n219_), .A2(new_n220_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT74), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n239_), .A2(new_n242_), .A3(KEYINPUT74), .A4(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT75), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n250_), .A3(new_n247_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT85), .B1(new_n259_), .B2(KEYINPUT1), .ZN(new_n260_));
  INV_X1    g059(.A(G155gat), .ZN(new_n261_));
  INV_X1    g060(.A(G162gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT86), .B1(new_n259_), .B2(KEYINPUT1), .ZN(new_n265_));
  OR3_X1    g064(.A1(new_n259_), .A2(KEYINPUT86), .A3(KEYINPUT1), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT84), .ZN(new_n269_));
  INV_X1    g068(.A(G141gat), .ZN(new_n270_));
  INV_X1    g069(.A(G148gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n269_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n269_), .A2(KEYINPUT87), .A3(new_n274_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n268_), .A2(new_n274_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n272_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT3), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n277_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G155gat), .B(G162gat), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT88), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT88), .B1(new_n284_), .B2(new_n285_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n273_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G113gat), .ZN(new_n291_));
  INV_X1    g090(.A(G120gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n273_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n284_), .A2(new_n285_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT88), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n296_), .B1(new_n299_), .B2(new_n286_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n293_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n295_), .A2(new_n301_), .A3(KEYINPUT4), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n300_), .A2(KEYINPUT4), .A3(new_n293_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n258_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n295_), .A2(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n258_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n257_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n257_), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n304_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT23), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n316_));
  MUX2_X1   g115(.A(new_n315_), .B(new_n316_), .S(KEYINPUT82), .Z(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(KEYINPUT24), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n320_), .A2(KEYINPUT24), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(G190gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT25), .B(G183gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n317_), .A2(new_n322_), .A3(new_n323_), .A4(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n315_), .B1(G183gat), .B2(G190gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G169gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n319_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n321_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G197gat), .B(G204gat), .Z(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(KEYINPUT91), .A3(KEYINPUT21), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n334_), .B(new_n335_), .C1(KEYINPUT21), .C2(new_n333_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n329_), .A2(KEYINPUT80), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n318_), .A2(KEYINPUT22), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n319_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n321_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT78), .B(G183gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n317_), .B1(G190gat), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n315_), .A2(new_n323_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n347_), .B2(KEYINPUT25), .ZN(new_n354_));
  INV_X1    g153(.A(new_n324_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n352_), .B(new_n322_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT92), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n338_), .B(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(KEYINPUT20), .B(new_n339_), .C1(new_n357_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n360_), .A2(KEYINPUT96), .A3(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT96), .B1(new_n360_), .B2(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n357_), .A2(new_n359_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n332_), .A2(new_n338_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT20), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n362_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT18), .B(G64gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G92gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n360_), .A2(new_n362_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n362_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n365_), .A2(KEYINPUT20), .A3(new_n377_), .A4(new_n366_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n374_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(KEYINPUT27), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383_));
  INV_X1    g182(.A(new_n379_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(new_n373_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n385_), .B2(new_n380_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G15gat), .B(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n293_), .B(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G71gat), .B(G99gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT31), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n357_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n349_), .A2(new_n356_), .A3(new_n394_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n392_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n399_), .A2(new_n400_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n391_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G22gat), .B(G50gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n289_), .B2(KEYINPUT29), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT29), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n300_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n232_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n418_), .B(new_n359_), .C1(new_n300_), .C2(new_n407_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n289_), .A2(KEYINPUT29), .B1(new_n337_), .B2(new_n336_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(new_n418_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n406_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n413_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425_));
  INV_X1    g224(.A(new_n422_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n411_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n424_), .B(KEYINPUT93), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n419_), .B(new_n430_), .C1(new_n420_), .C2(new_n418_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n423_), .A2(new_n424_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT94), .B1(new_n413_), .B2(new_n422_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n421_), .A2(new_n429_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n404_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n428_), .A2(new_n432_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n413_), .A2(new_n424_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n439_));
  AND4_X1   g238(.A1(new_n404_), .A2(new_n436_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n313_), .B(new_n387_), .C1(new_n437_), .C2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n311_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n379_), .B(new_n373_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n311_), .B(new_n446_), .C1(new_n304_), .C2(new_n308_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n302_), .A2(new_n303_), .A3(new_n258_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n306_), .A2(new_n307_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n257_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .A4(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n369_), .A2(KEYINPUT32), .A3(new_n373_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT32), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n384_), .B1(new_n453_), .B2(new_n374_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n452_), .B(new_n454_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n433_), .A2(new_n436_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n404_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n253_), .B1(new_n441_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G190gat), .B(G218gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G134gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(new_n262_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT36), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G232gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT68), .Z(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT34), .Z(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  INV_X1    g269(.A(G43gat), .ZN(new_n471_));
  INV_X1    g270(.A(G29gat), .ZN(new_n472_));
  INV_X1    g271(.A(G36gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G29gat), .A2(G36gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n471_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(G50gat), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(G50gat), .B1(new_n477_), .B2(new_n478_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n470_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G50gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n478_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n476_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n479_), .A3(KEYINPUT15), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT10), .B(G99gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT9), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G85gat), .A2(G92gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT9), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n499_), .A2(KEYINPUT64), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT64), .B1(new_n499_), .B2(new_n502_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n496_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n495_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n508_), .A2(new_n490_), .A3(new_n491_), .A4(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n497_), .A2(new_n498_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n510_), .A2(new_n511_), .A3(new_n516_), .A4(new_n512_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n505_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n487_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n480_), .A2(new_n481_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n520_), .A2(new_n505_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n521_));
  AOI211_X1 g320(.A(new_n465_), .B(new_n469_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n468_), .A2(KEYINPUT35), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n469_), .A2(new_n465_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n519_), .A2(new_n521_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n464_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n521_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT35), .A3(new_n468_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n463_), .A4(new_n525_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n460_), .B1(new_n527_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT69), .B1(new_n522_), .B2(new_n526_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n535_), .A3(new_n525_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n536_), .A3(new_n464_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT70), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n534_), .A2(new_n536_), .A3(new_n539_), .A4(new_n464_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n538_), .A2(new_n460_), .A3(new_n531_), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n533_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n459_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n520_), .A2(new_n229_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n487_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n547_), .B(new_n548_), .C1(new_n549_), .C2(new_n229_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n228_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n547_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G113gat), .B(G141gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(G169gat), .B(G197gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n550_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n505_), .A2(new_n515_), .A3(new_n214_), .A4(new_n517_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n515_), .A2(new_n517_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n490_), .B(new_n491_), .C1(new_n493_), .C2(G106gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n499_), .A2(new_n502_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT64), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n499_), .A2(KEYINPUT64), .A3(new_n502_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n241_), .B(new_n569_), .C1(new_n570_), .C2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n569_), .B1(new_n518_), .B2(new_n241_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n565_), .B(new_n568_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n241_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n566_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(G230gat), .A3(G233gat), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G204gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT5), .ZN(new_n587_));
  INV_X1    g386(.A(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n585_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT5), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(new_n591_), .A3(G176gat), .ZN(new_n592_));
  AOI21_X1  g391(.A(G176gat), .B1(new_n587_), .B2(new_n591_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n584_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(KEYINPUT67), .A3(new_n592_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT67), .ZN(new_n597_));
  INV_X1    g396(.A(new_n592_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n593_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(new_n584_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT13), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n546_), .A2(new_n564_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n313_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n223_), .A3(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT97), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(KEYINPUT97), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT38), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT98), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n441_), .A2(new_n458_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n538_), .A2(new_n540_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n531_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n602_), .A2(new_n564_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n612_), .A2(new_n248_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n313_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n606_), .A2(new_n621_), .A3(KEYINPUT38), .A4(new_n607_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n610_), .A2(new_n611_), .A3(new_n620_), .A4(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  INV_X1    g423(.A(new_n387_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n224_), .B1(new_n618_), .B2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT39), .Z(new_n627_));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n603_), .A2(new_n224_), .A3(new_n625_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n624_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(KEYINPUT40), .A3(new_n630_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n404_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n603_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT100), .Z(new_n640_));
  AOI21_X1  g439(.A(new_n637_), .B1(new_n618_), .B2(new_n638_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT41), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n457_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n618_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT101), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n603_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(new_n545_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n612_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(KEYINPUT102), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n545_), .B1(new_n441_), .B2(new_n458_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(KEYINPUT43), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n252_), .A2(new_n616_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n659_), .A2(KEYINPUT103), .A3(new_n660_), .A4(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n654_), .A2(KEYINPUT102), .A3(new_n652_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n656_), .B2(new_n657_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n661_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n660_), .A2(KEYINPUT103), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n651_), .B1(new_n670_), .B2(new_n313_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(KEYINPUT104), .A3(new_n604_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(G29gat), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n614_), .B1(new_n441_), .B2(new_n458_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(new_n661_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n472_), .A3(new_n604_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n473_), .A3(new_n625_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT45), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n387_), .B1(new_n662_), .B2(new_n668_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT105), .B(new_n679_), .C1(new_n680_), .C2(new_n473_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT106), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n680_), .B2(new_n473_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT105), .B1(new_n685_), .B2(new_n683_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n682_), .A2(new_n683_), .B1(new_n684_), .B2(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n675_), .A2(new_n471_), .A3(new_n638_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n404_), .B1(new_n662_), .B2(new_n668_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n471_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1330gat));
  AOI21_X1  g491(.A(G50gat), .B1(new_n675_), .B2(new_n645_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n670_), .A2(new_n483_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n645_), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n602_), .A2(new_n564_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n459_), .A2(new_n614_), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT107), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(G57gat), .A3(new_n604_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n546_), .A2(new_n696_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n202_), .B1(new_n700_), .B2(new_n313_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1332gat));
  AOI21_X1  g501(.A(new_n203_), .B1(new_n698_), .B2(new_n625_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT48), .Z(new_n704_));
  INV_X1    g503(.A(new_n700_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n203_), .A3(new_n625_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n698_), .B2(new_n638_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT49), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n705_), .A2(new_n708_), .A3(new_n638_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1334gat));
  INV_X1    g511(.A(G78gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n698_), .B2(new_n645_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT50), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n705_), .A2(new_n713_), .A3(new_n645_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1335gat));
  INV_X1    g516(.A(G85gat), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n253_), .A2(new_n696_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n674_), .A2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n721_), .B2(new_n313_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT108), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n655_), .A2(new_n658_), .A3(new_n719_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n313_), .A2(new_n718_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n724_), .B2(new_n725_), .ZN(G1336gat));
  NAND3_X1  g525(.A1(new_n724_), .A2(G92gat), .A3(new_n625_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n721_), .A2(new_n387_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(G92gat), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT109), .ZN(G1337gat));
  AOI21_X1  g529(.A(new_n507_), .B1(new_n724_), .B2(new_n638_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n721_), .A2(new_n493_), .A3(new_n404_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n724_), .A2(new_n645_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G106gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT52), .B(new_n495_), .C1(new_n724_), .C2(new_n645_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n645_), .A2(new_n495_), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n737_), .A2(new_n738_), .B1(new_n721_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g540(.A(new_n564_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n545_), .A2(new_n252_), .A3(new_n742_), .A4(new_n602_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT54), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n596_), .A2(new_n599_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT55), .B(new_n568_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(KEYINPUT110), .A2(G230gat), .A3(G233gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n748_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n580_), .B2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n745_), .B1(new_n753_), .B2(KEYINPUT56), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n580_), .A2(new_n751_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n748_), .A3(new_n747_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n566_), .A2(new_n567_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n569_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n581_), .A2(new_n759_), .ZN(new_n760_));
  AOI211_X1 g559(.A(new_n751_), .B(new_n758_), .C1(new_n760_), .C2(new_n577_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n600_), .B1(new_n761_), .B2(new_n750_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(KEYINPUT111), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n755_), .A3(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n564_), .A2(new_n595_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(KEYINPUT112), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT112), .B1(new_n766_), .B2(new_n767_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n553_), .B(new_n548_), .C1(new_n549_), .C2(new_n229_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n552_), .A2(new_n547_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n561_), .A3(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n563_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n601_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n768_), .A2(new_n769_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT57), .B1(new_n776_), .B2(new_n615_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n769_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n766_), .A2(KEYINPUT112), .A3(new_n767_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n774_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n614_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n595_), .A2(new_n773_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n783_), .A2(KEYINPUT113), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT113), .ZN(new_n785_));
  INV_X1    g584(.A(new_n755_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n753_), .A2(KEYINPUT56), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n784_), .B(new_n785_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT58), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n777_), .A2(new_n782_), .B1(new_n653_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n744_), .B1(new_n790_), .B2(new_n248_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n625_), .A2(new_n313_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(new_n437_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n564_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n777_), .A2(new_n782_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n653_), .A2(new_n789_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n253_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n790_), .B2(new_n252_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n744_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n793_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT59), .B1(new_n793_), .B2(new_n805_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT116), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n804_), .A2(new_n810_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n742_), .B(new_n797_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n795_), .B1(new_n812_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g612(.A(new_n292_), .B1(new_n602_), .B2(KEYINPUT60), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n794_), .B(new_n814_), .C1(KEYINPUT60), .C2(new_n292_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT117), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n602_), .B(new_n797_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n292_), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n794_), .B2(new_n252_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n248_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n797_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g621(.A(G134gat), .B1(new_n794_), .B2(new_n615_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n797_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n653_), .A2(G134gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(G1343gat));
  AND2_X1   g625(.A1(new_n791_), .A2(new_n440_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n792_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n742_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(new_n270_), .ZN(G1344gat));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n602_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(new_n271_), .ZN(G1345gat));
  NOR2_X1   g631(.A1(new_n828_), .A2(new_n253_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT61), .B(G155gat), .Z(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(G1346gat));
  NOR3_X1   g634(.A1(new_n828_), .A2(new_n262_), .A3(new_n545_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n827_), .A2(new_n615_), .A3(new_n792_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n262_), .B2(new_n837_), .ZN(G1347gat));
  NAND3_X1  g637(.A1(new_n625_), .A2(new_n313_), .A3(new_n638_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n742_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT118), .Z(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n645_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n318_), .B1(new_n804_), .B2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(KEYINPUT62), .Z(new_n844_));
  NOR2_X1   g643(.A1(new_n839_), .A2(new_n645_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n804_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n564_), .A2(new_n329_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n846_), .B2(new_n847_), .ZN(G1348gat));
  NAND2_X1  g647(.A1(new_n791_), .A2(new_n457_), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n849_), .A2(new_n319_), .A3(new_n602_), .A4(new_n839_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n602_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n804_), .A2(new_n851_), .A3(new_n845_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n319_), .ZN(G1349gat));
  NOR2_X1   g652(.A1(new_n820_), .A2(new_n325_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n804_), .A2(new_n845_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT119), .ZN(new_n856_));
  INV_X1    g655(.A(new_n347_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n839_), .A2(new_n253_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n849_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n804_), .A2(new_n860_), .A3(new_n845_), .A4(new_n854_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT120), .ZN(G1350gat));
  OAI21_X1  g662(.A(G190gat), .B1(new_n846_), .B2(new_n545_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n615_), .A2(new_n324_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT121), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n846_), .B2(new_n866_), .ZN(G1351gat));
  NAND3_X1  g666(.A1(new_n440_), .A2(KEYINPUT122), .A3(new_n313_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT122), .B1(new_n440_), .B2(new_n313_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n387_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n248_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n743_), .B(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n868_), .B(new_n870_), .C1(new_n871_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n791_), .A2(KEYINPUT123), .A3(new_n868_), .A4(new_n870_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n564_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT124), .B(G197gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1352gat));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n851_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n588_), .A2(KEYINPUT125), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1353gat));
  AOI21_X1  g683(.A(new_n820_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT126), .Z(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1354gat));
  INV_X1    g688(.A(G218gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n878_), .B2(new_n653_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n614_), .A2(G218gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT127), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n545_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n896_), .B(new_n897_), .C1(new_n890_), .C2(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n895_), .A2(new_n899_), .ZN(G1355gat));
endmodule


