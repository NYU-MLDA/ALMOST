//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G155gat), .B(G162gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G155gat), .ZN(new_n220_));
  INV_X1    g019(.A(G162gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G155gat), .A3(G162gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n221_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G141gat), .B(G148gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G127gat), .B(G134gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n229_), .A2(new_n234_), .A3(KEYINPUT92), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n217_), .A2(new_n218_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT92), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n236_), .A2(new_n237_), .B1(new_n233_), .B2(new_n232_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT4), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n236_), .A2(new_n234_), .A3(KEYINPUT4), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n208_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n234_), .B1(new_n229_), .B2(KEYINPUT92), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n230_), .B(new_n231_), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n208_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n207_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n247_), .B1(new_n252_), .B2(new_n240_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n246_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n208_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n255_), .A3(new_n206_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(new_n250_), .A3(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n253_), .A2(new_n255_), .A3(KEYINPUT97), .A4(new_n206_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G8gat), .B(G36gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT18), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT32), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT23), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT23), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(G183gat), .A3(G190gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n268_), .A3(KEYINPUT83), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n265_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n270_));
  NOR3_X1   g069(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n269_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT25), .B(G183gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(KEYINPUT24), .A3(new_n279_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n277_), .A2(KEYINPUT91), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT91), .B1(new_n277_), .B2(new_n280_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n274_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(G197gat), .A2(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT21), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G218gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G211gat), .ZN(new_n291_));
  INV_X1    g090(.A(G211gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G218gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n286_), .B(new_n289_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n293_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT87), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n266_), .A2(new_n268_), .ZN(new_n304_));
  OR2_X1    g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n283_), .A2(new_n303_), .A3(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n269_), .A2(new_n270_), .A3(new_n305_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n280_), .A2(KEYINPUT82), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT26), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT26), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n275_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n271_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n278_), .A2(new_n320_), .A3(KEYINPUT24), .A4(new_n279_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n313_), .A2(new_n318_), .A3(new_n319_), .A4(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n312_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n297_), .A2(new_n302_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n310_), .A2(KEYINPUT20), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT19), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(KEYINPUT96), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT96), .B1(new_n326_), .B2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n277_), .A2(new_n280_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT91), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n277_), .A2(KEYINPUT91), .A3(new_n280_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n273_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n309_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n324_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(KEYINPUT90), .B(KEYINPUT20), .C1(new_n323_), .C2(new_n324_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n303_), .A2(new_n312_), .A3(new_n322_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT90), .B1(new_n341_), .B2(KEYINPUT20), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n340_), .A2(new_n342_), .A3(new_n328_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n264_), .B1(new_n331_), .B2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n259_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n328_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n328_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n310_), .A2(KEYINPUT20), .A3(new_n348_), .A4(new_n325_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n349_), .A3(new_n264_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT95), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n263_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n263_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n253_), .A2(new_n255_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT33), .B1(new_n356_), .B2(new_n207_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n206_), .B1(new_n254_), .B2(new_n208_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n239_), .A2(new_n208_), .A3(new_n241_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n239_), .A2(KEYINPUT94), .A3(new_n208_), .A4(new_n241_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n364_), .B(new_n206_), .C1(new_n253_), .C2(new_n255_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n357_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n346_), .A2(new_n351_), .B1(new_n355_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n374_), .A3(new_n324_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n370_), .B2(new_n324_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n369_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n324_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n373_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n369_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G22gat), .B(G50gat), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n385_));
  NOR3_X1   g184(.A1(new_n229_), .A2(KEYINPUT29), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n236_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n384_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n236_), .A2(new_n388_), .A3(new_n387_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n383_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n378_), .A2(new_n382_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n378_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n381_), .B1(new_n380_), .B2(new_n375_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT88), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n399_), .A3(new_n382_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT86), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n394_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n390_), .A2(new_n393_), .A3(KEYINPUT86), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI211_X1 g203(.A(new_n368_), .B(new_n395_), .C1(new_n400_), .C2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n382_), .B1(new_n398_), .B2(KEYINPUT88), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n378_), .A2(new_n396_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n395_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT89), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n405_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT98), .B1(new_n367_), .B2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n357_), .A2(new_n363_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n354_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n365_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n413_), .A2(new_n352_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n343_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n258_), .B(new_n257_), .C1(new_n417_), .C2(new_n264_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n350_), .B(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT98), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n405_), .A2(new_n410_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT27), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n263_), .B(KEYINPUT99), .Z(new_n427_));
  NOR2_X1   g226(.A1(new_n417_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n352_), .A2(KEYINPUT27), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n411_), .A3(new_n259_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n412_), .A2(new_n424_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G227gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(G71gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G99gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n323_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(new_n234_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT84), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT30), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT31), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n439_), .B(new_n443_), .Z(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n433_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n431_), .A2(new_n423_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n259_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT75), .B(G8gat), .ZN(new_n452_));
  INV_X1    g251(.A(G1gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT14), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G1gat), .B(G8gat), .Z(new_n457_));
  OR2_X1    g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G29gat), .B(G36gat), .Z(new_n462_));
  XOR2_X1   g261(.A(G43gat), .B(G50gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT15), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G229gat), .A2(G233gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n464_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n471_), .A2(new_n467_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(new_n468_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G113gat), .B(G141gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT79), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G169gat), .B(G197gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n473_), .A2(KEYINPUT80), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n473_), .B2(KEYINPUT80), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G134gat), .B(G162gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(G190gat), .B(G218gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT36), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT73), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT74), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT70), .ZN(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n489_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT6), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G85gat), .ZN(new_n501_));
  INV_X1    g300(.A(G92gat), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT9), .ZN(new_n503_));
  XOR2_X1   g302(.A(G85gat), .B(G92gat), .Z(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(KEYINPUT9), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n495_), .A2(new_n500_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT65), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT65), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n510_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n500_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G99gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n489_), .A3(KEYINPUT66), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT66), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT67), .B(new_n504_), .C1(new_n512_), .C2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(new_n500_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n524_), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n504_), .A3(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n504_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT68), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT69), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n523_), .A2(new_n504_), .A3(new_n525_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n524_), .B1(new_n523_), .B2(new_n504_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n521_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n507_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n465_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n488_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n521_), .A2(new_n528_), .A3(new_n506_), .A4(new_n526_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n539_), .B(new_n544_), .C1(new_n545_), .C2(new_n470_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n533_), .A2(new_n464_), .A3(new_n506_), .A4(new_n521_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n539_), .B1(new_n548_), .B2(new_n544_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n534_), .B1(new_n533_), .B2(new_n521_), .ZN(new_n551_));
  AND4_X1   g350(.A1(new_n534_), .A2(new_n521_), .A3(new_n526_), .A4(new_n528_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n506_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(KEYINPUT70), .A3(new_n465_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n538_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n542_), .A2(new_n543_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n556_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n548_), .A2(new_n558_), .A3(new_n544_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n553_), .B2(new_n465_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n487_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n484_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT72), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n560_), .B(new_n566_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT37), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n557_), .A2(new_n561_), .A3(new_n565_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n560_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n569_), .B(new_n570_), .C1(new_n571_), .C2(new_n486_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G57gat), .B(G64gat), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT11), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT11), .ZN(new_n576_));
  XOR2_X1   g375(.A(G71gat), .B(G78gat), .Z(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n461_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT76), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(KEYINPUT76), .ZN(new_n585_));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n590_));
  OR4_X1    g389(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n589_), .B(KEYINPUT17), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT78), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n573_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n598_));
  INV_X1    g397(.A(new_n580_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT12), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n545_), .A2(new_n599_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT12), .B1(new_n545_), .B2(new_n599_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n553_), .A2(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n545_), .B(new_n599_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(G230gat), .A3(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT5), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n606_), .A2(new_n608_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n613_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n598_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(KEYINPUT13), .A3(new_n614_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n597_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n451_), .A2(new_n481_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT100), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n449_), .B1(new_n433_), .B2(new_n445_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n481_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n621_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n259_), .A2(G1gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n623_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT101), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n623_), .A2(new_n628_), .A3(new_n632_), .A4(new_n629_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(KEYINPUT38), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n259_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n569_), .B1(new_n571_), .B2(new_n486_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n624_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n620_), .A2(new_n625_), .A3(new_n595_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(KEYINPUT102), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT102), .B1(new_n638_), .B2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G1gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT38), .B1(new_n631_), .B2(new_n633_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT103), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n631_), .A2(new_n633_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n643_), .A4(new_n634_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n651_), .ZN(G1324gat));
  NAND3_X1  g451(.A1(new_n638_), .A2(new_n430_), .A3(new_n639_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n623_), .A2(new_n628_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n430_), .A2(new_n452_), .ZN(new_n658_));
  OAI22_X1  g457(.A1(new_n655_), .A2(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n659_), .B(new_n661_), .ZN(G1325gat));
  OR3_X1    g461(.A1(new_n622_), .A2(G15gat), .A3(new_n445_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n640_), .A2(new_n641_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n444_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n665_), .B2(G15gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n423_), .A2(KEYINPUT105), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n423_), .A2(KEYINPUT105), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n664_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n669_), .B1(new_n673_), .B2(G22gat), .ZN(new_n674_));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT42), .B(new_n675_), .C1(new_n664_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n672_), .A2(new_n675_), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n674_), .A2(new_n676_), .B1(new_n622_), .B2(new_n677_), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n637_), .A2(new_n595_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n620_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n626_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n635_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n624_), .B2(new_n573_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n573_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n259_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n430_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n421_), .A2(new_n423_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(KEYINPUT98), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n444_), .B1(new_n690_), .B2(new_n424_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n685_), .B(new_n686_), .C1(new_n691_), .C2(new_n449_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n684_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n620_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(new_n481_), .A3(new_n595_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n684_), .B2(new_n692_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n699_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n635_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n683_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  XNOR2_X1  g507(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n431_), .A2(G36gat), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n681_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n681_), .B2(new_n711_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n430_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI221_X1 g520(.A(new_n715_), .B1(KEYINPUT108), .B2(KEYINPUT46), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  INV_X1    g522(.A(G43gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n445_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n701_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n700_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n705_), .B(new_n725_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n681_), .B2(new_n445_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT47), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n732_), .A3(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n682_), .B2(new_n672_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n411_), .A2(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n706_), .B2(new_n736_), .ZN(G1331gat));
  NOR3_X1   g536(.A1(new_n694_), .A2(new_n481_), .A3(new_n595_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n638_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n638_), .A2(KEYINPUT110), .A3(new_n738_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n635_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G57gat), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n624_), .A2(new_n481_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n597_), .A2(new_n694_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n259_), .A2(G57gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n744_), .B1(new_n749_), .B2(new_n750_), .ZN(G1332gat));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n430_), .A3(new_n742_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(G64gat), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G64gat), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n431_), .A2(G64gat), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n754_), .A2(new_n755_), .B1(new_n749_), .B2(new_n756_), .ZN(G1333gat));
  NAND3_X1  g556(.A1(new_n741_), .A2(new_n444_), .A3(new_n742_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G71gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G71gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n444_), .A2(new_n435_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n760_), .A2(new_n761_), .B1(new_n749_), .B2(new_n762_), .ZN(G1334gat));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n747_), .A2(new_n764_), .A3(new_n672_), .A4(new_n748_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n741_), .A2(new_n672_), .A3(new_n742_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G78gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT112), .B(new_n765_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1335gat));
  NAND3_X1  g573(.A1(new_n620_), .A2(new_n625_), .A3(new_n595_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n684_), .B2(new_n692_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n259_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n679_), .A2(new_n694_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n747_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n635_), .A2(new_n501_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(G1336gat));
  OAI21_X1  g581(.A(G92gat), .B1(new_n777_), .B2(new_n431_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n430_), .A2(new_n502_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n780_), .B2(new_n784_), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n777_), .B2(new_n445_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n493_), .A2(new_n494_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n444_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n780_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI211_X1 g589(.A(new_n423_), .B(new_n775_), .C1(new_n684_), .C2(new_n692_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n489_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n776_), .A2(new_n411_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(G106gat), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n792_), .A2(new_n795_), .A3(KEYINPUT52), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT113), .B(new_n797_), .C1(new_n791_), .C2(new_n489_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n747_), .A2(new_n489_), .A3(new_n411_), .A4(new_n779_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT53), .B1(new_n796_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(new_n795_), .A3(KEYINPUT52), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n798_), .A3(new_n803_), .A4(new_n799_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT55), .B1(new_n605_), .B2(KEYINPUT114), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n530_), .A2(new_n535_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n600_), .B1(new_n809_), .B2(new_n506_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n603_), .A2(new_n602_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n603_), .A2(new_n602_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n807_), .B1(KEYINPUT55), .B2(new_n605_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n813_), .B(new_n815_), .C1(new_n536_), .C2(new_n600_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n612_), .A4(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n613_), .B1(new_n604_), .B2(new_n815_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n812_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  INV_X1    g621(.A(new_n812_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n816_), .A2(new_n612_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n819_), .A2(new_n821_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n473_), .A2(new_n478_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n468_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n466_), .A2(new_n467_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n471_), .B2(new_n467_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n477_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n614_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n826_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n568_), .A4(new_n572_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT58), .B1(new_n826_), .B2(new_n833_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT116), .B1(new_n573_), .B2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n834_), .A2(new_n835_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n825_), .A2(new_n817_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n481_), .A3(new_n614_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n832_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n847_), .B2(new_n636_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n595_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n694_), .A2(new_n573_), .A3(new_n625_), .A4(new_n596_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n852_), .A2(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n447_), .A2(new_n445_), .A3(new_n259_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT117), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n806_), .B1(new_n860_), .B2(new_n625_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n861_), .A2(KEYINPUT118), .ZN(new_n862_));
  INV_X1    g661(.A(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT119), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n859_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n850_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n843_), .A2(new_n849_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(KEYINPUT120), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n843_), .A2(new_n872_), .A3(new_n849_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n596_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n868_), .B1(new_n874_), .B2(new_n855_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n855_), .B1(new_n595_), .B2(new_n851_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n876_), .B2(new_n863_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n875_), .A2(G113gat), .A3(new_n481_), .A4(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n861_), .A2(KEYINPUT118), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n862_), .A2(new_n878_), .A3(new_n879_), .ZN(G1340gat));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n573_), .A2(new_n839_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n841_), .B1(new_n883_), .B2(new_n837_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n848_), .B1(new_n884_), .B2(new_n840_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n850_), .B1(new_n885_), .B2(new_n872_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n873_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n595_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n882_), .B1(new_n888_), .B2(new_n856_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n863_), .B1(new_n852_), .B2(new_n856_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n620_), .B1(new_n890_), .B2(new_n867_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n881_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n875_), .A2(KEYINPUT122), .A3(new_n620_), .A4(new_n877_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(G120gat), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT121), .B1(new_n895_), .B2(G120gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(G120gat), .B1(new_n620_), .B2(new_n895_), .ZN(new_n897_));
  MUX2_X1   g696(.A(new_n896_), .B(KEYINPUT121), .S(new_n897_), .Z(new_n898_));
  NAND2_X1  g697(.A1(new_n890_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n899_), .ZN(G1341gat));
  INV_X1    g699(.A(G127gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n595_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n870_), .A2(KEYINPUT120), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n850_), .A3(new_n873_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n855_), .B1(new_n904_), .B2(new_n595_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n877_), .B(new_n902_), .C1(new_n905_), .C2(new_n882_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n901_), .B1(new_n860_), .B2(new_n595_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(KEYINPUT123), .A3(new_n907_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1342gat));
  NAND3_X1  g711(.A1(new_n875_), .A2(new_n686_), .A3(new_n877_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G134gat), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n636_), .A2(G134gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n860_), .B2(new_n915_), .ZN(G1343gat));
  NOR4_X1   g715(.A1(new_n423_), .A2(new_n430_), .A3(new_n444_), .A4(new_n259_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n876_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n481_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n620_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g722(.A1(new_n857_), .A2(new_n917_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n924_), .B2(new_n595_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n919_), .A2(new_n926_), .A3(new_n596_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT61), .B(G155gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1346gat));
  OAI21_X1  g729(.A(G162gat), .B1(new_n924_), .B2(new_n573_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n919_), .A2(new_n221_), .A3(new_n637_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n431_), .A2(new_n448_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n672_), .A2(new_n935_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n481_), .B(new_n936_), .C1(new_n874_), .C2(new_n855_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n937_), .A2(new_n938_), .A3(G169gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n937_), .B2(G169gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n936_), .B1(new_n874_), .B2(new_n855_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT22), .B(G169gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n481_), .A2(new_n942_), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n943_), .B(KEYINPUT125), .Z(new_n944_));
  OAI22_X1  g743(.A1(new_n939_), .A2(new_n940_), .B1(new_n941_), .B2(new_n944_), .ZN(G1348gat));
  INV_X1    g744(.A(new_n941_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G176gat), .B1(new_n946_), .B2(new_n620_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n876_), .A2(new_n411_), .A3(new_n935_), .ZN(new_n948_));
  INV_X1    g747(.A(G176gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n694_), .A2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n948_), .B2(new_n950_), .ZN(G1349gat));
  AOI21_X1  g750(.A(G183gat), .B1(new_n948_), .B2(new_n596_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n595_), .A2(new_n275_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n946_), .B2(new_n953_), .ZN(G1350gat));
  OAI21_X1  g753(.A(G190gat), .B1(new_n941_), .B2(new_n573_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n637_), .A2(new_n276_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n941_), .B2(new_n956_), .ZN(G1351gat));
  NOR3_X1   g756(.A1(new_n431_), .A2(new_n687_), .A3(new_n444_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n876_), .A2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n481_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n620_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  NAND4_X1  g765(.A1(new_n960_), .A2(new_n596_), .A3(new_n965_), .A4(new_n966_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  AND2_X1   g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n857_), .A2(new_n958_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n595_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n967_), .B1(new_n971_), .B2(new_n965_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n969_), .B1(new_n972_), .B2(KEYINPUT126), .ZN(G1354gat));
  NOR2_X1   g772(.A1(new_n970_), .A2(new_n573_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n637_), .A2(new_n290_), .ZN(new_n975_));
  OAI22_X1  g774(.A1(new_n974_), .A2(new_n290_), .B1(new_n970_), .B2(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(KEYINPUT127), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978_));
  OAI221_X1 g777(.A(new_n978_), .B1(new_n970_), .B2(new_n975_), .C1(new_n974_), .C2(new_n290_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n977_), .A2(new_n979_), .ZN(G1355gat));
endmodule


