//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT79), .ZN(new_n206_));
  INV_X1    g005(.A(new_n204_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n203_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT79), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n206_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT31), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G71gat), .B(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G43gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n219_), .A2(new_n221_), .B1(KEYINPUT24), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT25), .B(G183gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT26), .B(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n225_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n233_), .B2(new_n232_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n238_));
  OAI21_X1  g037(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n239_));
  OR3_X1    g038(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n242_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n244_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n217_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT77), .B(G15gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n244_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n216_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT80), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n251_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n213_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n254_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n251_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n261_), .A2(KEYINPUT80), .A3(new_n255_), .A4(new_n212_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G197gat), .B(G204gat), .Z(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT21), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n274_), .B(new_n276_), .Z(new_n277_));
  AND2_X1   g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT82), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(G155gat), .B2(G162gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT2), .ZN(new_n286_));
  OR2_X1    g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT3), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(KEYINPUT3), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n288_), .B(new_n289_), .C1(new_n285_), .C2(KEYINPUT2), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n282_), .B1(new_n286_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT1), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n287_), .B(new_n283_), .C1(new_n281_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT29), .ZN(new_n296_));
  INV_X1    g095(.A(G228gat), .ZN(new_n297_));
  INV_X1    g096(.A(G233gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n278_), .A2(new_n296_), .A3(KEYINPUT87), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n272_), .A2(new_n277_), .A3(new_n300_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n302_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n295_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n278_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n301_), .A2(new_n306_), .B1(new_n309_), .B2(new_n299_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n307_), .A2(new_n304_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G22gat), .B(G50gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT28), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n319_), .B(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n316_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT89), .B1(new_n310_), .B2(new_n312_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n322_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n324_), .A2(KEYINPUT90), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n315_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n318_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT90), .B1(new_n324_), .B2(new_n325_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n314_), .A4(new_n313_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n232_), .B1(KEYINPUT91), .B2(new_n225_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(KEYINPUT91), .B2(new_n225_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n241_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n278_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n272_), .A2(new_n277_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(new_n241_), .A3(new_n235_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n278_), .A2(new_n242_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n337_), .A2(new_n241_), .A3(new_n334_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n341_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT20), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT18), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(new_n351_), .A3(new_n346_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(KEYINPUT92), .A3(new_n354_), .ZN(new_n355_));
  OR3_X1    g154(.A1(new_n347_), .A2(KEYINPUT92), .A3(new_n352_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(KEYINPUT27), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n343_), .A2(KEYINPUT20), .A3(new_n344_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n341_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n336_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n351_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(new_n359_), .A2(KEYINPUT94), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n206_), .A2(new_n210_), .A3(new_n295_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n307_), .A2(new_n205_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT4), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n367_), .A2(new_n369_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n373_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n373_), .B2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT94), .B1(new_n359_), .B2(new_n363_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n358_), .A2(new_n364_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n331_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n355_), .A2(new_n356_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n381_), .A2(KEYINPUT33), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(KEYINPUT33), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n378_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n368_), .A2(new_n372_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n390_), .B(KEYINPUT93), .C1(new_n391_), .C2(new_n370_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n370_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n327_), .A2(new_n330_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n361_), .A2(new_n362_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n351_), .A2(KEYINPUT32), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI221_X1 g200(.A(new_n401_), .B1(new_n347_), .B2(new_n400_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n258_), .A2(KEYINPUT81), .A3(new_n262_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n265_), .A2(new_n385_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT95), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n258_), .A2(KEYINPUT81), .A3(new_n262_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT81), .B1(new_n258_), .B2(new_n262_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n403_), .A4(new_n385_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n358_), .A2(new_n364_), .A3(new_n383_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n331_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n263_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n364_), .A2(new_n383_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(new_n398_), .A3(KEYINPUT96), .A4(new_n358_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n406_), .A2(new_n411_), .B1(new_n418_), .B2(new_n382_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G29gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G43gat), .B(G50gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT15), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT71), .B(G15gat), .ZN(new_n424_));
  INV_X1    g223(.A(G22gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT72), .B(G1gat), .Z(new_n427_));
  INV_X1    g226(.A(G8gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT14), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G8gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n423_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT75), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n431_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n422_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G229gat), .A2(G233gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  OR3_X1    g241(.A1(new_n438_), .A2(KEYINPUT74), .A3(new_n422_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n438_), .A2(new_n422_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT74), .A3(new_n439_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n443_), .A2(new_n446_), .A3(G229gat), .A4(G233gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G141gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G169gat), .B(G197gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n442_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n419_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G230gat), .A2(G233gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT64), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(KEYINPUT66), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n464_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n463_), .A2(new_n465_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G85gat), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n473_), .A2(new_n464_), .A3(KEYINPUT9), .A4(new_n461_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  AND2_X1   g274(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR4_X1   g279(.A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT65), .A4(G106gat), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n470_), .B(new_n474_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n473_), .A2(new_n461_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n467_), .A2(new_n469_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT8), .B(new_n483_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT8), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n479_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n468_), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n484_), .B(new_n493_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n483_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n490_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n482_), .B1(new_n489_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  INV_X1    g302(.A(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G57gat), .ZN(new_n505_));
  INV_X1    g304(.A(G57gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G64gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n502_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n499_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n482_), .B(new_n511_), .C1(new_n489_), .C2(new_n498_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(KEYINPUT12), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n499_), .A2(new_n516_), .A3(new_n512_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n460_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n519_), .A3(new_n514_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n467_), .A2(new_n469_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n493_), .A2(new_n484_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n497_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT8), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n496_), .A2(new_n490_), .A3(new_n497_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n511_), .B1(new_n526_), .B2(new_n482_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n459_), .B1(new_n527_), .B2(KEYINPUT67), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n518_), .B1(new_n520_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n534_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n535_), .A2(KEYINPUT13), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT13), .B1(new_n535_), .B2(new_n536_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n420_), .B(new_n421_), .Z(new_n540_));
  NAND2_X1  g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT34), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n499_), .A2(new_n540_), .B1(KEYINPUT35), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n423_), .A2(new_n499_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546_));
  INV_X1    g345(.A(new_n542_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n544_), .B(new_n545_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n546_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n545_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n543_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT68), .B(KEYINPUT36), .Z(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT37), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n548_), .A2(new_n551_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n548_), .A2(new_n551_), .A3(KEYINPUT69), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n557_), .ZN(new_n567_));
  OAI211_X1 g366(.A(KEYINPUT70), .B(new_n561_), .C1(new_n567_), .C2(KEYINPUT37), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n511_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n438_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT17), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n571_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT73), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n566_), .A2(new_n583_), .A3(new_n584_), .A4(new_n557_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n539_), .A2(new_n568_), .A3(new_n582_), .A4(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n457_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n382_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n427_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591_));
  OAI22_X1  g390(.A1(new_n588_), .A2(new_n590_), .B1(KEYINPUT98), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT98), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(new_n567_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n419_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n539_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n581_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n456_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(KEYINPUT97), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(KEYINPUT97), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n603_), .B2(new_n382_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n594_), .A2(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(KEYINPUT40), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n413_), .A3(new_n599_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n428_), .B1(new_n608_), .B2(KEYINPUT100), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(KEYINPUT39), .A3(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n457_), .A2(new_n428_), .A3(new_n413_), .A4(new_n587_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT99), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT39), .B1(new_n609_), .B2(new_n611_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n606_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n618_), .A2(KEYINPUT40), .A3(new_n612_), .A4(new_n614_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1325gat));
  OR3_X1    g419(.A1(new_n588_), .A2(G15gat), .A3(new_n409_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n409_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n623_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT41), .B1(new_n623_), .B2(G15gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(G1326gat));
  XNOR2_X1  g425(.A(new_n331_), .B(KEYINPUT101), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT42), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n629_), .A2(new_n630_), .A3(G22gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n629_), .B2(G22gat), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n425_), .ZN(new_n633_));
  OAI22_X1  g432(.A1(new_n631_), .A2(new_n632_), .B1(new_n588_), .B2(new_n633_), .ZN(G1327gat));
  XOR2_X1   g433(.A(new_n581_), .B(KEYINPUT73), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n595_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT103), .ZN(new_n637_));
  NOR4_X1   g436(.A1(new_n419_), .A2(new_n456_), .A3(new_n597_), .A4(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(G29gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n589_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n406_), .A2(new_n411_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n418_), .A2(new_n382_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT37), .B(new_n558_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n561_), .A2(KEYINPUT70), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n585_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n582_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n597_), .A2(new_n456_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(KEYINPUT43), .A3(new_n646_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n650_), .A4(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n646_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n419_), .B2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n651_), .A2(new_n654_), .A3(new_n650_), .A4(new_n635_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n652_), .A2(new_n657_), .A3(new_n589_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(KEYINPUT102), .ZN(new_n659_));
  OAI21_X1  g458(.A(G29gat), .B1(new_n658_), .B2(KEYINPUT102), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n640_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n657_), .A3(new_n413_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  INV_X1    g462(.A(G36gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n638_), .A2(new_n664_), .A3(new_n413_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n663_), .A2(new_n666_), .A3(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  NAND3_X1  g470(.A1(new_n652_), .A2(new_n657_), .A3(new_n415_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G43gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n638_), .A2(new_n215_), .A3(new_n622_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT47), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(KEYINPUT47), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1330gat));
  INV_X1    g478(.A(G50gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n638_), .A2(new_n680_), .A3(new_n628_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n652_), .A2(new_n657_), .A3(new_n331_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n682_), .A2(KEYINPUT104), .ZN(new_n683_));
  OAI21_X1  g482(.A(G50gat), .B1(new_n682_), .B2(KEYINPUT104), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(G1331gat));
  NOR2_X1   g484(.A1(new_n419_), .A2(new_n455_), .ZN(new_n686_));
  AND4_X1   g485(.A1(new_n597_), .A2(new_n686_), .A3(new_n582_), .A4(new_n653_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n506_), .A3(new_n589_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n539_), .A2(new_n455_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n643_), .A2(new_n567_), .A3(new_n582_), .A4(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G57gat), .B1(new_n690_), .B2(new_n382_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1332gat));
  NAND2_X1  g491(.A1(new_n413_), .A2(new_n504_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT105), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n413_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G64gat), .B1(new_n690_), .B2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT106), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n690_), .B2(new_n409_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n687_), .A2(new_n704_), .A3(new_n622_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1334gat));
  OAI21_X1  g505(.A(G78gat), .B1(new_n690_), .B2(new_n627_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT50), .ZN(new_n708_));
  INV_X1    g507(.A(G78gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n687_), .A2(new_n709_), .A3(new_n628_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n637_), .A2(new_n539_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n686_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n471_), .A3(new_n589_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n649_), .A2(KEYINPUT107), .A3(new_n651_), .A4(new_n689_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n651_), .A2(new_n654_), .A3(new_n635_), .A4(new_n689_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n382_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n719_), .B2(new_n471_), .ZN(G1336gat));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n472_), .A3(new_n413_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n696_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n472_), .ZN(G1337gat));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n415_), .A3(new_n478_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT108), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n409_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n492_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT51), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n725_), .C1(new_n726_), .C2(new_n492_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1338gat));
  NAND4_X1  g530(.A1(new_n686_), .A2(new_n479_), .A3(new_n331_), .A4(new_n712_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  OAI21_X1  g534(.A(G106gat), .B1(new_n716_), .B2(new_n398_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n735_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT53), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n736_), .A2(new_n735_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n738_), .A4(new_n734_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT59), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n418_), .A2(new_n589_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n586_), .A2(new_n455_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  NOR4_X1   g549(.A1(new_n586_), .A2(new_n750_), .A3(KEYINPUT54), .A4(new_n455_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT110), .B1(new_n747_), .B2(new_n748_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n567_), .A2(KEYINPUT57), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n455_), .A2(new_n536_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n759_), .B(new_n760_), .C1(new_n518_), .C2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n514_), .A2(KEYINPUT12), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n527_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n517_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n459_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT114), .B1(new_n766_), .B2(KEYINPUT111), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT55), .B1(new_n518_), .B2(new_n759_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT112), .B1(new_n764_), .B2(new_n765_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n515_), .A2(new_n772_), .A3(new_n517_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n460_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT113), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n515_), .A2(new_n517_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n459_), .B1(new_n776_), .B2(KEYINPUT112), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n773_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n533_), .B1(new_n770_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n769_), .A2(new_n775_), .A3(new_n779_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n533_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n758_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n440_), .B1(new_n438_), .B2(new_n422_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n451_), .B1(new_n437_), .B2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n446_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT115), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n535_), .A2(new_n536_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n437_), .A2(new_n787_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n452_), .A4(new_n789_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n791_), .A2(new_n792_), .A3(new_n454_), .A4(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n757_), .B1(new_n786_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n536_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n802_));
  AND4_X1   g601(.A1(new_n778_), .A2(new_n771_), .A3(new_n460_), .A4(new_n773_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n778_), .B1(new_n777_), .B2(new_n773_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI211_X1 g604(.A(new_n782_), .B(new_n534_), .C1(new_n805_), .C2(new_n769_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n533_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n796_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT117), .A3(new_n757_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n800_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n567_), .B1(new_n786_), .B2(new_n797_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n795_), .A2(new_n454_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n794_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n801_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n653_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n817_), .B(KEYINPUT58), .C1(new_n806_), .C2(new_n807_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n812_), .A2(new_n814_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n582_), .B1(new_n811_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n755_), .B1(new_n823_), .B2(KEYINPUT119), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n825_), .B(new_n582_), .C1(new_n811_), .C2(new_n822_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n745_), .B(new_n746_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n811_), .A2(new_n822_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n598_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n829_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n755_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(new_n746_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n834_), .B2(new_n745_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n456_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n837_), .A3(new_n455_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1340gat));
  OAI21_X1  g638(.A(G120gat), .B1(new_n835_), .B2(new_n539_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n539_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n834_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n834_), .B2(new_n582_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n835_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n581_), .A2(G127gat), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT120), .Z(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n846_), .B2(new_n848_), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n835_), .B2(new_n653_), .ZN(new_n850_));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n834_), .A2(new_n851_), .A3(new_n595_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n622_), .A2(new_n398_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n413_), .A2(new_n382_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n833_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n455_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n856_), .A2(new_n539_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT121), .B(G148gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n856_), .A2(new_n635_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT61), .B(G155gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  INV_X1    g664(.A(G162gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n857_), .B2(new_n646_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n856_), .A2(G162gat), .A3(new_n567_), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n867_), .A2(KEYINPUT122), .A3(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT122), .B1(new_n867_), .B2(new_n868_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1347gat));
  NOR3_X1   g670(.A1(new_n409_), .A2(new_n589_), .A3(new_n696_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n455_), .A3(new_n627_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n753_), .A2(new_n749_), .A3(new_n751_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT117), .B1(new_n809_), .B2(new_n757_), .ZN(new_n875_));
  AOI211_X1 g674(.A(new_n799_), .B(new_n756_), .C1(new_n808_), .C2(new_n796_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n791_), .A2(new_n454_), .A3(new_n536_), .A4(new_n795_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n646_), .B1(new_n879_), .B2(KEYINPUT58), .ZN(new_n880_));
  INV_X1    g679(.A(new_n821_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n595_), .B1(new_n808_), .B2(new_n796_), .ZN(new_n882_));
  OAI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n882_), .B2(new_n813_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n635_), .B1(new_n877_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n874_), .B1(new_n884_), .B2(new_n825_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n823_), .A2(KEYINPUT119), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n873_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT22), .B(G169gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  OAI21_X1  g689(.A(G169gat), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  AOI211_X1 g690(.A(KEYINPUT123), .B(new_n873_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n891_), .A2(KEYINPUT62), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  INV_X1    g693(.A(new_n873_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n222_), .B1(new_n896_), .B2(KEYINPUT123), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n887_), .A2(new_n890_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n889_), .B1(new_n893_), .B2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n889_), .C1(new_n893_), .C2(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1348gat));
  NAND2_X1  g703(.A1(new_n872_), .A2(new_n627_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n906_), .B2(new_n597_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n833_), .A2(new_n398_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n872_), .A2(G176gat), .A3(new_n597_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n907_), .B1(new_n910_), .B2(new_n912_), .ZN(G1349gat));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n582_), .A3(new_n872_), .ZN(new_n914_));
  INV_X1    g713(.A(G183gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n598_), .A2(new_n226_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n914_), .A2(new_n915_), .B1(new_n906_), .B2(new_n916_), .ZN(G1350gat));
  NAND2_X1  g716(.A1(new_n906_), .A2(new_n646_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G190gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n906_), .A2(new_n227_), .A3(new_n595_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n696_), .A2(new_n589_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n833_), .A2(new_n854_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT126), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n833_), .A2(new_n925_), .A3(new_n854_), .A4(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n927_), .A2(G197gat), .A3(new_n455_), .ZN(new_n928_));
  AOI21_X1  g727(.A(G197gat), .B1(new_n927_), .B2(new_n455_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1352gat));
  AOI21_X1  g729(.A(new_n539_), .B1(new_n924_), .B2(new_n926_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT127), .B(G204gat), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1353gat));
  XNOR2_X1  g732(.A(KEYINPUT63), .B(G211gat), .ZN(new_n934_));
  AOI211_X1 g733(.A(new_n598_), .B(new_n934_), .C1(new_n924_), .C2(new_n926_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n927_), .A2(new_n581_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n927_), .A2(new_n939_), .A3(new_n595_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n653_), .B1(new_n924_), .B2(new_n926_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(new_n941_), .ZN(G1355gat));
endmodule


