//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT34), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT70), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n218_), .A3(KEYINPUT64), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n214_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n216_), .A2(new_n218_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT66), .B(new_n212_), .C1(new_n231_), .C2(new_n229_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n219_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT66), .B1(new_n234_), .B2(new_n212_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n230_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237_));
  OR2_X1    g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n226_), .A3(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n210_), .A2(KEYINPUT9), .A3(new_n211_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n237_), .B1(new_n223_), .B2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n245_), .A2(KEYINPUT65), .A3(new_n222_), .A4(new_n221_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT15), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n207_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n212_), .B1(new_n231_), .B2(new_n229_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT8), .A3(new_n232_), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n258_), .A2(new_n230_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n259_), .B2(new_n251_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n236_), .A2(new_n254_), .A3(new_n247_), .A4(new_n251_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n253_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n204_), .A2(new_n205_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n236_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT69), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n264_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n253_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G190gat), .B(G218gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT71), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G134gat), .B(G162gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT36), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT72), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n265_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n274_), .B(KEYINPUT36), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n268_), .A2(new_n269_), .A3(new_n253_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n269_), .B1(new_n268_), .B2(new_n253_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n279_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT73), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n202_), .B(KEYINPUT37), .C1(new_n283_), .C2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT37), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n284_), .A2(new_n285_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n286_), .A2(KEYINPUT73), .B1(new_n290_), .B2(new_n277_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n281_), .A2(new_n282_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n286_), .A2(new_n278_), .A3(new_n289_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT74), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT75), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n298_), .B(new_n288_), .C1(new_n293_), .C2(new_n295_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G1gat), .ZN(new_n301_));
  INV_X1    g100(.A(G8gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT14), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n303_), .A2(KEYINPUT76), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(KEYINPUT76), .ZN(new_n305_));
  XOR2_X1   g104(.A(G15gat), .B(G22gat), .Z(new_n306_));
  NOR3_X1   g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G8gat), .Z(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G64gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT11), .ZN(new_n313_));
  XOR2_X1   g112(.A(G71gat), .B(G78gat), .Z(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n314_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(KEYINPUT11), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n315_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n311_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT17), .ZN(new_n324_));
  XOR2_X1   g123(.A(G127gat), .B(G155gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G183gat), .B(G211gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n323_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(KEYINPUT17), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G230gat), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n259_), .A2(new_n320_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n248_), .A2(new_n319_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT12), .ZN(new_n338_));
  OR3_X1    g137(.A1(new_n259_), .A2(KEYINPUT12), .A3(new_n320_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI211_X1 g139(.A(new_n333_), .B(new_n334_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G120gat), .B(G148gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT5), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G176gat), .B(G204gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT67), .B1(new_n342_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n342_), .B2(new_n347_), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT67), .B(new_n346_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT13), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT68), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n300_), .A2(new_n332_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G15gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G71gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G99gat), .ZN(new_n366_));
  INV_X1    g165(.A(G71gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n364_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n225_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT23), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G183gat), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G169gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(G176gat), .B1(new_n383_), .B2(KEYINPUT22), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT22), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n385_), .A3(G169gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n380_), .A2(new_n381_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT26), .B1(new_n375_), .B2(KEYINPUT80), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n374_), .A2(KEYINPUT25), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n395_));
  NOR2_X1   g194(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n396_));
  OAI21_X1  g195(.A(G183gat), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT79), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(G183gat), .C1(new_n395_), .C2(new_n396_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n394_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n378_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n377_), .A2(KEYINPUT23), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n381_), .A2(KEYINPUT24), .ZN(new_n406_));
  INV_X1    g205(.A(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(G176gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n404_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n388_), .B1(new_n401_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n388_), .B(KEYINPUT30), .C1(new_n401_), .C2(new_n411_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n370_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n370_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT83), .B(G43gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n414_), .A2(new_n415_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(new_n416_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n361_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n420_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(KEYINPUT84), .ZN(new_n428_));
  INV_X1    g227(.A(G134gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G127gat), .ZN(new_n430_));
  INV_X1    g229(.A(G127gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G134gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G120gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G113gat), .ZN(new_n435_));
  INV_X1    g234(.A(G113gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G120gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n430_), .A2(new_n432_), .A3(new_n435_), .A4(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT31), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n425_), .A2(new_n428_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n361_), .B(new_n444_), .C1(new_n421_), .C2(new_n424_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447_));
  INV_X1    g246(.A(G141gat), .ZN(new_n448_));
  INV_X1    g247(.A(G148gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G141gat), .A2(G148gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT2), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n450_), .A2(new_n453_), .A3(new_n454_), .A4(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT1), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n465_), .A3(new_n458_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n467_), .A2(new_n451_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n460_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n439_), .A2(new_n440_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT99), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n441_), .A2(new_n460_), .A3(new_n469_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(KEYINPUT99), .A3(new_n471_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT4), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT100), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G225gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n472_), .B2(KEYINPUT4), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n479_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT100), .B1(new_n486_), .B2(new_n482_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G29gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G85gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT0), .B(G57gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  AOI21_X1  g290(.A(new_n481_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n484_), .A2(new_n487_), .A3(new_n491_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n482_), .B1(new_n477_), .B2(KEYINPUT4), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n496_), .B2(new_n479_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n491_), .B1(new_n497_), .B2(new_n487_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT101), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n484_), .A2(new_n487_), .A3(new_n493_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n491_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT101), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n494_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n446_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT18), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G197gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT88), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G197gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n513_), .A3(G204gat), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n511_), .A2(new_n513_), .A3(KEYINPUT90), .A4(G204gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n510_), .B2(G204gat), .ZN(new_n520_));
  INV_X1    g319(.A(G204gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G211gat), .B(G218gat), .Z(new_n525_));
  NAND3_X1  g324(.A1(new_n511_), .A2(new_n513_), .A3(new_n521_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(G197gat), .B2(G204gat), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n516_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n525_), .A2(KEYINPUT21), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT20), .B1(new_n533_), .B2(new_n412_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n385_), .A2(G169gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n407_), .A2(KEYINPUT22), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n535_), .A2(new_n536_), .A3(KEYINPUT96), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT96), .B1(new_n535_), .B2(new_n536_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n408_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT81), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n377_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT23), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n403_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n376_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n381_), .B(KEYINPUT95), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n539_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT25), .B(G183gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT26), .B(G190gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n410_), .A2(new_n550_), .A3(new_n379_), .A4(new_n373_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n529_), .A2(new_n532_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n553_));
  AND2_X1   g352(.A1(G226gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT94), .Z(new_n556_));
  NOR3_X1   g355(.A1(new_n534_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n533_), .B2(new_n412_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n524_), .A2(new_n528_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n555_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n509_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT102), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n556_), .B1(new_n534_), .B2(new_n552_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n509_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n555_), .A3(new_n561_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT97), .B(new_n556_), .C1(new_n534_), .C2(new_n552_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT102), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n572_), .B(new_n509_), .C1(new_n557_), .C2(new_n562_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n564_), .A2(new_n571_), .A3(KEYINPUT27), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT103), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(KEYINPUT27), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT103), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n571_), .A4(new_n564_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n570_), .A2(new_n569_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n411_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n398_), .A2(new_n400_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n394_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n560_), .A2(new_n584_), .A3(new_n388_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n547_), .A2(new_n551_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n533_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n587_), .A3(KEYINPUT20), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT97), .B1(new_n588_), .B2(new_n556_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n509_), .B1(new_n579_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n571_), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n592_));
  AOI22_X1  g391(.A1(new_n575_), .A2(new_n578_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G78gat), .B(G106gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT87), .B1(new_n470_), .B2(KEYINPUT29), .ZN(new_n596_));
  NAND2_X1  g395(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(G233gat), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n470_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT91), .B1(new_n460_), .B2(new_n469_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT29), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n560_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n600_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n533_), .B2(new_n596_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n595_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n533_), .A2(new_n596_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n600_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n596_), .A2(new_n602_), .B1(new_n604_), .B2(KEYINPUT29), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n611_), .B(new_n594_), .C1(new_n612_), .C2(new_n560_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n611_), .B1(new_n612_), .B2(new_n560_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT92), .B1(new_n615_), .B2(new_n595_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n470_), .A2(KEYINPUT29), .ZN(new_n617_));
  XOR2_X1   g416(.A(G22gat), .B(G50gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT28), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n617_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n614_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n609_), .A2(new_n613_), .A3(KEYINPUT92), .A4(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n505_), .A2(new_n593_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n575_), .A2(new_n578_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n591_), .A2(new_n592_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n609_), .A2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n631_), .A2(new_n620_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n623_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n502_), .A2(new_n503_), .A3(new_n494_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n503_), .B1(new_n502_), .B2(new_n494_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n629_), .B(new_n634_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n627_), .B1(new_n628_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n575_), .A2(new_n578_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n624_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(KEYINPUT105), .A4(new_n629_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n591_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n472_), .A2(KEYINPUT4), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n486_), .A2(new_n481_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n480_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n645_), .A2(new_n491_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n494_), .A2(KEYINPUT33), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n497_), .A2(new_n649_), .A3(new_n491_), .A4(new_n487_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n590_), .A2(KEYINPUT98), .A3(new_n571_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n643_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n568_), .A2(KEYINPUT32), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n567_), .A2(new_n569_), .A3(new_n570_), .A4(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n557_), .A2(new_n562_), .ZN(new_n656_));
  OAI221_X1 g455(.A(new_n655_), .B1(new_n656_), .B2(new_n654_), .C1(new_n495_), .C2(new_n498_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n624_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n638_), .A2(new_n641_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n626_), .B1(new_n660_), .B2(new_n446_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n311_), .A2(new_n252_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n309_), .A2(new_n251_), .A3(new_n310_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(G229gat), .A2(G233gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n311_), .B(new_n251_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n664_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(G113gat), .B(G141gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G169gat), .B(G197gat), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n668_), .B(new_n669_), .Z(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n667_), .B(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n661_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n360_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n499_), .A2(new_n504_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(new_n301_), .A3(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT38), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n286_), .A2(new_n278_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n661_), .A2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT107), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n357_), .B2(new_n673_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT106), .B(new_n672_), .C1(new_n353_), .C2(new_n356_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n332_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n684_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G1gat), .B1(new_n689_), .B2(new_n677_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n680_), .A2(new_n690_), .ZN(G1324gat));
  INV_X1    g490(.A(new_n593_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n676_), .A2(new_n302_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT39), .ZN(new_n694_));
  INV_X1    g493(.A(new_n689_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n692_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(G8gat), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT39), .B(new_n302_), .C1(new_n695_), .C2(new_n692_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g499(.A(G15gat), .B1(new_n689_), .B2(new_n446_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT41), .Z(new_n702_));
  INV_X1    g501(.A(new_n446_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n676_), .A2(new_n363_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1326gat));
  OAI21_X1  g504(.A(G22gat), .B1(new_n689_), .B2(new_n624_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT42), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n624_), .A2(G22gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n675_), .B2(new_n708_), .ZN(G1327gat));
  INV_X1    g508(.A(new_n332_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n682_), .ZN(new_n711_));
  NOR4_X1   g510(.A1(new_n661_), .A2(new_n673_), .A3(new_n357_), .A4(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G29gat), .B1(new_n712_), .B2(new_n678_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n299_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT37), .B1(new_n283_), .B2(new_n287_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n294_), .A2(KEYINPUT74), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n298_), .B1(new_n717_), .B2(new_n288_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n714_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n639_), .A2(new_n640_), .A3(new_n629_), .ZN(new_n721_));
  AOI22_X1  g520(.A1(new_n721_), .A2(new_n627_), .B1(new_n658_), .B2(new_n624_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n703_), .B1(new_n722_), .B2(new_n641_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n719_), .B(new_n720_), .C1(new_n723_), .C2(new_n626_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n661_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n727_), .A2(KEYINPUT109), .A3(new_n720_), .A4(new_n719_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n661_), .B2(new_n300_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n686_), .A2(new_n710_), .A3(new_n687_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT108), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n686_), .A2(new_n733_), .A3(new_n710_), .A4(new_n687_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n730_), .A2(KEYINPUT44), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT44), .B1(new_n730_), .B2(new_n735_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n678_), .A2(G29gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n713_), .B1(new_n738_), .B2(new_n739_), .ZN(G1328gat));
  NOR2_X1   g539(.A1(new_n593_), .A2(G36gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n712_), .A2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT45), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT45), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n661_), .A2(new_n300_), .A3(KEYINPUT43), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n729_), .B1(new_n747_), .B2(KEYINPUT109), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n724_), .A2(new_n725_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n735_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n730_), .A2(KEYINPUT44), .A3(new_n735_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n692_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n746_), .B1(new_n754_), .B2(G36gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT111), .B1(new_n755_), .B2(KEYINPUT46), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n755_), .B2(KEYINPUT110), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n759_), .B(new_n746_), .C1(new_n754_), .C2(G36gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n736_), .A2(new_n737_), .A3(new_n593_), .ZN(new_n762_));
  INV_X1    g561(.A(G36gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n745_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n759_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n755_), .A2(KEYINPUT110), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(KEYINPUT111), .A3(new_n757_), .A4(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n761_), .A2(new_n767_), .ZN(G1329gat));
  AOI21_X1  g567(.A(G43gat), .B1(new_n712_), .B2(new_n703_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT113), .Z(new_n770_));
  AND2_X1   g569(.A1(new_n703_), .A2(G43gat), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n738_), .A2(KEYINPUT112), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT112), .B1(new_n738_), .B2(new_n771_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g574(.A(G50gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n712_), .A2(new_n776_), .A3(new_n634_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n738_), .A2(KEYINPUT114), .A3(new_n634_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G50gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT114), .B1(new_n738_), .B2(new_n634_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(G1331gat));
  NOR2_X1   g580(.A1(new_n661_), .A2(new_n672_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n719_), .A2(new_n710_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n357_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT115), .ZN(new_n785_));
  AOI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n678_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT116), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n358_), .A2(new_n710_), .A3(new_n672_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n684_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n678_), .A2(G57gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(G1332gat));
  OAI21_X1  g591(.A(G64gat), .B1(new_n789_), .B2(new_n593_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n785_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n593_), .A2(G64gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(G1333gat));
  OAI21_X1  g597(.A(G71gat), .B1(new_n789_), .B2(new_n446_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT49), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n785_), .A2(new_n367_), .A3(new_n703_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1334gat));
  OAI21_X1  g601(.A(G78gat), .B1(new_n789_), .B2(new_n624_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n624_), .A2(G78gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n796_), .B2(new_n806_), .ZN(G1335gat));
  NOR2_X1   g606(.A1(new_n358_), .A2(new_n711_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n782_), .A2(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n809_), .A2(G85gat), .A3(new_n677_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n748_), .A2(new_n749_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n357_), .A2(new_n710_), .A3(new_n673_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n678_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n814_), .B2(G85gat), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT119), .Z(G1336gat));
  INV_X1    g615(.A(new_n809_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n209_), .A3(new_n692_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n811_), .A2(new_n593_), .A3(new_n812_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n209_), .ZN(G1337gat));
  NAND4_X1  g619(.A1(new_n817_), .A2(new_n703_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n811_), .A2(new_n446_), .A3(new_n812_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n225_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n813_), .A2(new_n634_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G106gat), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n809_), .A2(G106gat), .A3(new_n624_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  AOI211_X1 g631(.A(KEYINPUT120), .B(new_n226_), .C1(new_n813_), .C2(new_n634_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n827_), .A2(new_n833_), .A3(new_n828_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT53), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n830_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n827_), .A2(new_n828_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n836_), .B(new_n837_), .C1(new_n838_), .C2(new_n833_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(new_n839_), .ZN(G1339gat));
  NOR4_X1   g639(.A1(new_n692_), .A2(new_n677_), .A3(new_n634_), .A4(new_n446_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n667_), .A2(new_n671_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n664_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n662_), .A2(new_n663_), .A3(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n844_), .B(new_n671_), .C1(new_n666_), .C2(new_n843_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n842_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n349_), .A2(new_n350_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n340_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n338_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n340_), .A2(new_n848_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n346_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT56), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n342_), .A2(new_n347_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n851_), .A2(new_n856_), .A3(new_n346_), .A4(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n847_), .B1(new_n858_), .B2(new_n673_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n681_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n854_), .A2(new_n857_), .A3(new_n855_), .A4(new_n846_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT58), .Z(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n300_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n710_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n783_), .A2(new_n867_), .A3(new_n673_), .A4(new_n358_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n359_), .B2(new_n672_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n866_), .A2(new_n870_), .A3(KEYINPUT121), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT121), .B1(new_n866_), .B2(new_n870_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n841_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n436_), .A3(new_n672_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n841_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n870_), .B2(new_n866_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n873_), .B2(KEYINPUT59), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n879_), .A2(new_n672_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT122), .B(new_n875_), .C1(new_n880_), .C2(new_n436_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n436_), .B1(new_n879_), .B2(new_n672_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n875_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n885_), .ZN(G1340gat));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n887_));
  AOI21_X1  g686(.A(G120gat), .B1(new_n357_), .B2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT123), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n887_), .B2(G120gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n874_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n879_), .A2(new_n357_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n434_), .B2(new_n894_), .ZN(G1341gat));
  AOI21_X1  g694(.A(G127gat), .B1(new_n874_), .B2(new_n332_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n896_), .A2(KEYINPUT125), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(KEYINPUT125), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n710_), .A2(new_n431_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n898_), .B1(new_n879_), .B2(new_n899_), .ZN(G1342gat));
  NAND3_X1  g699(.A1(new_n874_), .A2(new_n429_), .A3(new_n682_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n879_), .A2(new_n719_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n429_), .ZN(G1343gat));
  OR2_X1    g702(.A1(new_n871_), .A2(new_n872_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n703_), .A2(new_n624_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n692_), .A2(new_n677_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n448_), .A3(new_n672_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G141gat), .B1(new_n908_), .B2(new_n673_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1344gat));
  NAND3_X1  g711(.A1(new_n909_), .A2(new_n449_), .A3(new_n357_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G148gat), .B1(new_n908_), .B2(new_n358_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1345gat));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n909_), .A2(new_n332_), .A3(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n908_), .B2(new_n710_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1346gat));
  OAI21_X1  g719(.A(G162gat), .B1(new_n908_), .B2(new_n300_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n681_), .A2(G162gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n908_), .B2(new_n922_), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n593_), .A2(new_n678_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n703_), .ZN(new_n925_));
  AOI211_X1 g724(.A(new_n634_), .B(new_n925_), .C1(new_n870_), .C2(new_n866_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927_), .B2(new_n673_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(KEYINPUT62), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n928_), .A2(KEYINPUT62), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n926_), .B(new_n672_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n926_), .B2(new_n357_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n904_), .A2(new_n624_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n358_), .A2(new_n408_), .A3(new_n925_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(G1349gat));
  NOR2_X1   g735(.A1(new_n925_), .A2(new_n710_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G183gat), .B1(new_n934_), .B2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n634_), .B1(new_n866_), .B2(new_n870_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n925_), .A2(new_n548_), .A3(new_n710_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n927_), .B2(new_n300_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n926_), .A2(new_n549_), .A3(new_n682_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n904_), .A2(new_n905_), .A3(new_n924_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n946_), .B(new_n672_), .C1(KEYINPUT126), .C2(G197gat), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT126), .B(G197gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(new_n945_), .B2(new_n673_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1352gat));
  NOR2_X1   g749(.A1(new_n945_), .A2(new_n358_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(new_n521_), .ZN(G1353gat));
  NOR2_X1   g751(.A1(new_n945_), .A2(new_n710_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AND2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n956_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n946_), .B2(new_n682_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n719_), .A2(G218gat), .ZN(new_n959_));
  XOR2_X1   g758(.A(new_n959_), .B(KEYINPUT127), .Z(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n946_), .B2(new_n960_), .ZN(G1355gat));
endmodule


