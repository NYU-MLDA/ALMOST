//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT9), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT10), .B(G99gat), .ZN(new_n210_));
  OAI221_X1 g009(.A(new_n209_), .B1(KEYINPUT9), .B2(new_n208_), .C1(new_n210_), .C2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT66), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n211_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT67), .A3(new_n223_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n216_), .A3(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n207_), .A2(new_n208_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n224_), .A2(new_n225_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n218_), .A2(new_n235_), .A3(new_n219_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n221_), .B1(new_n234_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n242_));
  XOR2_X1   g041(.A(G71gat), .B(G78gat), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n237_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n232_), .A2(new_n237_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT66), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT66), .B1(new_n213_), .B2(new_n215_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n252_), .B2(new_n235_), .ZN(new_n253_));
  OAI22_X1  g052(.A1(new_n248_), .A2(new_n253_), .B1(new_n220_), .B2(new_n211_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n246_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n247_), .A2(KEYINPUT12), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n258_), .A3(new_n255_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n204_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n204_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n247_), .B2(new_n256_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT5), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(KEYINPUT68), .Z(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT13), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT13), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G232gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT34), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n281_), .B1(new_n254_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT15), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n285_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT15), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT71), .B1(new_n239_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(KEYINPUT15), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n254_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n287_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n279_), .A2(new_n280_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n276_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n239_), .A2(new_n289_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n254_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n294_), .B1(new_n254_), .B2(new_n295_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT72), .A3(new_n298_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n301_), .B(new_n299_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n293_), .A2(new_n296_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n310_), .A2(KEYINPUT74), .A3(new_n299_), .A4(new_n301_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G190gat), .B(G218gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G134gat), .B(G162gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT36), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT73), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n306_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT37), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n300_), .A2(new_n305_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n315_), .B(KEYINPUT36), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n319_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n306_), .A2(new_n312_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n323_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(KEYINPUT75), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n326_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n325_), .B1(new_n331_), .B2(KEYINPUT37), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G127gat), .B(G155gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT16), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G183gat), .B(G211gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G15gat), .B(G22gat), .ZN(new_n338_));
  INV_X1    g137(.A(G1gat), .ZN(new_n339_));
  INV_X1    g138(.A(G8gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT14), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G8gat), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G231gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(new_n246_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n337_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT17), .B1(new_n349_), .B2(new_n337_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(KEYINPUT17), .B(new_n337_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n332_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n275_), .A2(KEYINPUT77), .A3(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358_));
  INV_X1    g157(.A(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(G15gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n360_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT25), .B(G183gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT26), .B(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n365_), .A2(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n370_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n371_));
  AND2_X1   g170(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n372_));
  NOR2_X1   g171(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT84), .B1(new_n370_), .B2(KEYINPUT23), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n368_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT24), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G176gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(KEYINPUT85), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(G183gat), .B(G190gat), .C1(new_n372_), .C2(new_n373_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n370_), .A2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n380_), .A2(new_n391_), .A3(KEYINPUT30), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(KEYINPUT86), .A3(new_n395_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n364_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n364_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G127gat), .B(G134gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G113gat), .B(G120gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n403_), .A2(new_n404_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n400_), .A2(new_n402_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n409_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G141gat), .B(G148gat), .Z(new_n414_));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G155gat), .A3(G162gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT88), .ZN(new_n417_));
  INV_X1    g216(.A(G155gat), .ZN(new_n418_));
  INV_X1    g217(.A(G162gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(KEYINPUT87), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT1), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(G155gat), .B2(G162gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n414_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT91), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT2), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(G141gat), .A3(G148gat), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n428_), .A2(new_n430_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  AND2_X1   g235(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT90), .B(new_n436_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n435_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n420_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT92), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT92), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n420_), .A2(new_n424_), .A3(new_n446_), .A4(new_n421_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n426_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT29), .ZN(new_n450_));
  INV_X1    g249(.A(G204gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT95), .B1(new_n451_), .B2(G197gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  INV_X1    g252(.A(G197gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(G204gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(G197gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT21), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(new_n454_), .B2(G204gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT21), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n454_), .A2(G204gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G211gat), .B(G218gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n460_), .A2(new_n461_), .B1(new_n454_), .B2(G204gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n466_), .A2(new_n463_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G228gat), .A2(G233gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n450_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n435_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n478_), .B2(new_n426_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n466_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n468_), .B2(new_n463_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n481_), .A2(new_n458_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n475_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(new_n483_), .A3(KEYINPUT98), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G78gat), .B(G106gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT97), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n474_), .A2(new_n483_), .A3(KEYINPUT98), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(new_n449_), .B2(KEYINPUT29), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n478_), .A2(KEYINPUT93), .A3(new_n476_), .A4(new_n426_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G22gat), .B(G50gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n492_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n474_), .A2(new_n483_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT98), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n490_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n487_), .A2(new_n499_), .A3(new_n502_), .A4(new_n489_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G226gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT19), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n472_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n376_), .A2(new_n389_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n384_), .A2(KEYINPUT22), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n382_), .A2(G169gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n381_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(new_n378_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n386_), .A2(new_n388_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(new_n379_), .A3(new_n369_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n515_), .A2(new_n517_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n508_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT100), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G8gat), .B(G36gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n520_), .B(KEYINPUT100), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G64gat), .B(G92gat), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n482_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n392_), .A2(new_n472_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n508_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT20), .A4(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n519_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT105), .ZN(new_n539_));
  INV_X1    g338(.A(new_n533_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT20), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n369_), .A2(new_n379_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n542_), .A2(new_n516_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n543_), .B2(new_n482_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n536_), .B1(new_n544_), .B2(new_n535_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n509_), .A2(new_n518_), .A3(new_n508_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n540_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT105), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n519_), .A2(new_n533_), .A3(new_n548_), .A4(new_n537_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n539_), .A2(new_n547_), .A3(KEYINPUT27), .A4(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT27), .ZN(new_n551_));
  INV_X1    g350(.A(new_n538_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n533_), .B1(new_n519_), .B2(new_n537_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n449_), .A2(new_n407_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n407_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n478_), .A2(new_n557_), .A3(new_n426_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(KEYINPUT4), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G225gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT101), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n478_), .B2(new_n426_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT4), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n556_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G29gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G57gat), .B(G85gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n567_), .A3(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR4_X1   g376(.A1(new_n413_), .A2(new_n506_), .A3(new_n555_), .A4(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n555_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n567_), .A2(new_n573_), .ZN(new_n583_));
  AOI211_X1 g382(.A(new_n582_), .B(KEYINPUT33), .C1(new_n583_), .C2(new_n566_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT103), .B1(new_n576_), .B2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(KEYINPUT33), .A3(new_n566_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n553_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n556_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n559_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n560_), .B1(new_n556_), .B2(KEYINPUT4), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n574_), .B(new_n590_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n588_), .A2(new_n589_), .A3(new_n593_), .A4(new_n538_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n519_), .A2(new_n596_), .A3(new_n537_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n531_), .A2(KEYINPUT32), .A3(new_n532_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n546_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT20), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n508_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n598_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n519_), .A2(new_n537_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n587_), .A2(new_n595_), .B1(new_n577_), .B2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n581_), .B1(new_n607_), .B2(new_n506_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n578_), .B1(new_n608_), .B2(new_n413_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n346_), .A2(new_n286_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n289_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT78), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT78), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n346_), .A2(new_n615_), .A3(new_n286_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n288_), .A2(new_n346_), .A3(new_n291_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n613_), .A3(new_n611_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(KEYINPUT79), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT80), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT81), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT79), .B1(new_n617_), .B2(new_n619_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT82), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n617_), .A2(new_n619_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT79), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT82), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n620_), .A4(new_n625_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n609_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n357_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT77), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n275_), .A2(new_n356_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n339_), .A3(new_n577_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n609_), .A2(new_n331_), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n355_), .B(new_n636_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n577_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n643_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n644_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  NAND3_X1  g450(.A1(new_n641_), .A2(new_n340_), .A3(new_n555_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n555_), .A3(new_n646_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(G8gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G8gat), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n652_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n652_), .A2(new_n658_), .A3(KEYINPUT40), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647_), .B2(new_n413_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT107), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n641_), .A2(new_n362_), .A3(new_n412_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n506_), .B(KEYINPUT108), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n641_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G22gat), .B1(new_n647_), .B2(new_n673_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT42), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(G29gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n413_), .A2(new_n577_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n506_), .A2(new_n555_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n577_), .A2(new_n606_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n559_), .A2(new_n565_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n567_), .A2(new_n573_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n585_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n582_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n576_), .A2(KEYINPUT103), .A3(new_n585_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n683_), .B1(new_n689_), .B2(new_n594_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n506_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n690_), .A2(new_n691_), .B1(new_n580_), .B2(new_n579_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT109), .B(new_n682_), .C1(new_n692_), .C2(new_n412_), .ZN(new_n693_));
  AND2_X1   g492(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n693_), .B(new_n332_), .C1(new_n609_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n320_), .A2(new_n324_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n322_), .B1(new_n321_), .B2(KEYINPUT75), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n306_), .A2(KEYINPUT75), .A3(new_n312_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n319_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT37), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n696_), .B1(new_n609_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n273_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n355_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n636_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n695_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT110), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n708_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n709_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n679_), .B1(new_n714_), .B2(new_n577_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n331_), .A2(new_n355_), .ZN(new_n716_));
  NOR4_X1   g515(.A1(new_n609_), .A2(new_n704_), .A3(new_n716_), .A4(new_n636_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n718_), .A2(G29gat), .A3(new_n648_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT111), .B1(new_n715_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n709_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n713_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n712_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(new_n648_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726_));
  INV_X1    g525(.A(new_n719_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n714_), .B2(new_n555_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n555_), .A2(new_n731_), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n718_), .A2(KEYINPUT45), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT45), .B1(new_n718_), .B2(new_n733_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n730_), .B1(new_n732_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G36gat), .B1(new_n724_), .B2(new_n580_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(KEYINPUT46), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1329gat));
  NOR2_X1   g540(.A1(new_n413_), .A2(new_n359_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n721_), .B(new_n742_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n359_), .B1(new_n718_), .B2(new_n413_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g545(.A(G50gat), .B1(new_n717_), .B2(new_n674_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n506_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n714_), .B2(new_n748_), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n609_), .A2(new_n635_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n356_), .A3(new_n704_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n648_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n752_), .B2(new_n751_), .ZN(new_n754_));
  INV_X1    g553(.A(G57gat), .ZN(new_n755_));
  INV_X1    g554(.A(new_n275_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n355_), .A2(new_n635_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n645_), .A3(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n648_), .A2(new_n755_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n754_), .A2(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1332gat));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761_));
  INV_X1    g560(.A(G64gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n758_), .B2(new_n555_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n763_), .A2(new_n764_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n761_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n767_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT48), .A3(new_n765_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n751_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n762_), .A3(new_n555_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n770_), .A3(new_n772_), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n758_), .B2(new_n412_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT49), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n412_), .A2(new_n774_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT114), .Z(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n751_), .B2(new_n778_), .ZN(G1334gat));
  INV_X1    g578(.A(G78gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n758_), .B2(new_n674_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT50), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n771_), .A2(new_n780_), .A3(new_n674_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1335gat));
  NOR2_X1   g583(.A1(new_n275_), .A2(new_n716_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n750_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n205_), .A3(new_n577_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n704_), .A2(new_n355_), .A3(new_n636_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n695_), .A2(new_n703_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT115), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(KEYINPUT115), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n577_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n788_), .B1(new_n796_), .B2(new_n205_), .ZN(G1336gat));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n555_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G92gat), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n786_), .A2(G92gat), .A3(new_n580_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n206_), .B1(new_n794_), .B2(new_n555_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT116), .B1(new_n804_), .B2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1337gat));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT51), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(KEYINPUT51), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT118), .Z(new_n811_));
  INV_X1    g610(.A(new_n789_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n790_), .A2(KEYINPUT115), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n412_), .B(new_n812_), .C1(new_n813_), .C2(new_n791_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(G99gat), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n786_), .A2(new_n210_), .A3(new_n413_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n809_), .B(new_n811_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n811_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n814_), .B2(G99gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n808_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n812_), .A2(new_n695_), .A3(new_n506_), .A4(new_n703_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n822_), .A2(new_n823_), .A3(G106gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n822_), .B2(G106gat), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n691_), .A2(G106gat), .ZN(new_n826_));
  OAI22_X1  g625(.A1(new_n824_), .A2(new_n825_), .B1(new_n786_), .B2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g627(.A1(new_n681_), .A2(new_n577_), .A3(new_n412_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n257_), .A2(new_n259_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n261_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n257_), .A2(new_n204_), .A3(new_n259_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n269_), .B1(new_n260_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n635_), .A2(new_n268_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n611_), .A2(new_n614_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n624_), .B1(new_n842_), .B2(new_n618_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n612_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n629_), .A2(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n840_), .A2(new_n841_), .B1(new_n270_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT57), .B1(new_n847_), .B2(new_n331_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n839_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n835_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n841_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n270_), .A2(new_n846_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n700_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n268_), .A2(new_n846_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(KEYINPUT58), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n332_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n856_), .A2(new_n864_), .A3(new_n861_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n355_), .A3(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n702_), .A2(new_n273_), .A3(new_n757_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT54), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n636_), .B(new_n829_), .C1(new_n866_), .C2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT120), .B1(new_n869_), .B2(G113gat), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871_));
  INV_X1    g670(.A(G113gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n858_), .B(new_n873_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n848_), .A2(new_n855_), .B1(new_n874_), .B2(new_n332_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n355_), .B1(new_n875_), .B2(new_n864_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n865_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n868_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n829_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n871_), .B(new_n872_), .C1(new_n880_), .C2(new_n636_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n705_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT121), .B1(new_n875_), .B2(new_n705_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n868_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n880_), .A2(KEYINPUT59), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n636_), .A2(new_n872_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n870_), .A2(new_n881_), .B1(new_n888_), .B2(new_n889_), .ZN(G1340gat));
  AOI21_X1  g689(.A(new_n829_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n273_), .B2(KEYINPUT60), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n893_), .C1(KEYINPUT60), .C2(new_n892_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n886_), .A2(new_n887_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n895_), .B(new_n756_), .C1(new_n891_), .C2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n894_), .B1(new_n898_), .B2(new_n892_), .ZN(G1341gat));
  INV_X1    g698(.A(G127gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n891_), .A2(new_n900_), .A3(new_n705_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n895_), .B(new_n705_), .C1(new_n891_), .C2(new_n896_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n903_), .B2(new_n900_), .ZN(G1342gat));
  INV_X1    g703(.A(G134gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n891_), .A2(new_n905_), .A3(new_n331_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n895_), .B(new_n332_), .C1(new_n891_), .C2(new_n896_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n908_), .B2(new_n905_), .ZN(G1343gat));
  NOR4_X1   g708(.A1(new_n691_), .A2(new_n648_), .A3(new_n555_), .A4(new_n412_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n878_), .A2(new_n635_), .A3(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g711(.A1(new_n878_), .A2(new_n756_), .A3(new_n910_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g713(.A1(new_n878_), .A2(new_n910_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n355_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT61), .B(G155gat), .Z(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1346gat));
  NOR3_X1   g717(.A1(new_n915_), .A2(new_n419_), .A3(new_n702_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n878_), .A2(new_n331_), .A3(new_n910_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(G162gat), .ZN(new_n922_));
  OAI211_X1 g721(.A(KEYINPUT122), .B(new_n419_), .C1(new_n915_), .C2(new_n700_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n919_), .B1(new_n922_), .B2(new_n923_), .ZN(G1347gat));
  NAND2_X1  g723(.A1(new_n680_), .A2(new_n555_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n674_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n886_), .A2(new_n635_), .A3(new_n926_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n384_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(KEYINPUT124), .A3(new_n928_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n886_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n926_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n936_), .A2(new_n511_), .A3(new_n512_), .A4(new_n635_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n927_), .B(new_n931_), .C1(new_n930_), .C2(new_n929_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n933_), .A2(new_n937_), .A3(new_n938_), .ZN(G1348gat));
  NAND2_X1  g738(.A1(new_n936_), .A2(new_n704_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n506_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n275_), .A2(new_n381_), .A3(new_n925_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n940_), .A2(new_n381_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  NOR4_X1   g742(.A1(new_n934_), .A2(new_n355_), .A3(new_n365_), .A4(new_n935_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n925_), .A2(new_n355_), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n878_), .A2(new_n691_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G183gat), .B1(new_n946_), .B2(KEYINPUT125), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n941_), .A2(new_n945_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n944_), .B1(new_n947_), .B2(new_n950_), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n936_), .A2(new_n331_), .A3(new_n366_), .ZN(new_n952_));
  INV_X1    g751(.A(G190gat), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n934_), .A2(new_n702_), .A3(new_n935_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n952_), .B1(new_n953_), .B2(new_n954_), .ZN(G1351gat));
  NAND3_X1  g754(.A1(new_n413_), .A2(new_n506_), .A3(new_n648_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n957_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n958_), .A2(new_n959_), .A3(new_n580_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n878_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n636_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(new_n454_), .ZN(G1352gat));
  NOR2_X1   g762(.A1(new_n961_), .A2(new_n275_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(new_n451_), .ZN(G1353gat));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  AND2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  NOR4_X1   g766(.A1(new_n961_), .A2(new_n355_), .A3(new_n966_), .A4(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n961_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n705_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n968_), .B1(new_n970_), .B2(new_n966_), .ZN(G1354gat));
  XNOR2_X1  g770(.A(KEYINPUT127), .B(G218gat), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n961_), .A2(new_n702_), .A3(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n969_), .A2(new_n331_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n974_), .B2(new_n972_), .ZN(G1355gat));
endmodule


