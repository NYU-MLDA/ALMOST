//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_;
  XNOR2_X1  g000(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G230gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  OAI22_X1  g009(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(new_n221_), .A3(new_n219_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT64), .B(G85gat), .ZN(new_n226_));
  INV_X1    g025(.A(G92gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n218_), .ZN(new_n230_));
  OR2_X1    g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n214_), .A3(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n229_), .A2(new_n210_), .A3(new_n230_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n225_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G64gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G57gat), .ZN(new_n237_));
  INV_X1    g036(.A(G57gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G64gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n239_), .A3(KEYINPUT11), .ZN(new_n243_));
  INV_X1    g042(.A(G78gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G71gat), .ZN(new_n245_));
  INV_X1    g044(.A(G71gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G78gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n242_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n250_), .A2(KEYINPUT11), .A3(new_n245_), .A4(new_n247_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT67), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(new_n248_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n254_), .B(new_n251_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n235_), .A2(KEYINPUT68), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260_));
  INV_X1    g059(.A(new_n257_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n254_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n234_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n260_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n235_), .A2(new_n258_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n205_), .B(new_n259_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n249_), .A2(KEYINPUT12), .A3(new_n251_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n216_), .A2(new_n221_), .A3(new_n219_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n221_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n234_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n230_), .A2(new_n210_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n278_), .A2(KEYINPUT69), .A3(new_n233_), .A4(new_n229_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n272_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n263_), .A2(new_n265_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n270_), .A2(new_n204_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G120gat), .B(G148gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(G176gat), .B(G204gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n268_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n268_), .B2(new_n283_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n203_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n268_), .A2(new_n283_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n268_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT71), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n291_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT34), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT35), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G43gat), .B(G50gat), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n309_), .B(new_n234_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n302_), .A2(KEYINPUT35), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n307_), .A2(KEYINPUT15), .A3(new_n308_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT15), .B1(new_n307_), .B2(new_n308_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n275_), .B2(new_n280_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n304_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT15), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n309_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n307_), .A2(KEYINPUT15), .A3(new_n308_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n277_), .A2(new_n279_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(new_n225_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n310_), .A2(new_n312_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n303_), .B(KEYINPUT74), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G190gat), .B(G218gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G134gat), .B(G162gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n320_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n319_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n338_), .B2(new_n304_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n332_), .B(KEYINPUT36), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n335_), .B(KEYINPUT75), .C1(new_n339_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT37), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G155gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT16), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G183gat), .B(G211gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT17), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(KEYINPUT77), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(KEYINPUT17), .ZN(new_n351_));
  AND2_X1   g150(.A1(G15gat), .A2(G22gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G15gat), .A2(G22gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT14), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(G1gat), .B2(G8gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G15gat), .B(G22gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359_));
  INV_X1    g158(.A(G1gat), .ZN(new_n360_));
  INV_X1    g159(.A(G8gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT14), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(G1gat), .B(G8gat), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n357_), .A2(new_n365_), .A3(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(G231gat), .A3(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G231gat), .A2(G233gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n367_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n252_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n370_), .A2(new_n251_), .A3(new_n249_), .A4(new_n373_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n349_), .A2(new_n254_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n348_), .ZN(new_n380_));
  AOI211_X1 g179(.A(new_n350_), .B(new_n351_), .C1(new_n377_), .C2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(new_n378_), .A3(new_n376_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n320_), .A2(new_n329_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n340_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(KEYINPUT75), .A3(KEYINPUT37), .A4(new_n335_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n300_), .A2(new_n344_), .A3(new_n383_), .A4(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT101), .ZN(new_n388_));
  INV_X1    g187(.A(G169gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT22), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT22), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G169gat), .ZN(new_n392_));
  INV_X1    g191(.A(G176gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT82), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT22), .B(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n395_), .A2(new_n398_), .B1(G169gat), .B2(G176gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT23), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT23), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(G183gat), .A3(G190gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n403_), .A3(KEYINPUT83), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n400_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n405_));
  INV_X1    g204(.A(G183gat), .ZN(new_n406_));
  INV_X1    g205(.A(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(KEYINPUT25), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT25), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G183gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(KEYINPUT26), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT26), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G190gat), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .A4(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(KEYINPUT24), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT24), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n416_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n400_), .B2(KEYINPUT23), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n402_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n401_), .A3(new_n426_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n399_), .A2(new_n409_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT84), .B(G15gat), .Z(new_n429_));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n428_), .B(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n428_), .A2(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n428_), .A2(new_n431_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G71gat), .B(G99gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G43gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT30), .ZN(new_n442_));
  XOR2_X1   g241(.A(G127gat), .B(G134gat), .Z(new_n443_));
  INV_X1    g242(.A(G120gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G113gat), .ZN(new_n445_));
  INV_X1    g244(.A(G113gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(G120gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT85), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n448_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G127gat), .B(G134gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G113gat), .B(G120gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n449_), .B1(new_n454_), .B2(KEYINPUT85), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n442_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n439_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT0), .B(G57gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G141gat), .ZN(new_n463_));
  INV_X1    g262(.A(G148gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n465_), .A2(KEYINPUT3), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT87), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT87), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(new_n474_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n468_), .A2(new_n473_), .A3(new_n476_), .A4(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G155gat), .B(G162gat), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n465_), .A2(new_n467_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT1), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n481_), .A2(new_n486_), .A3(new_n454_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n443_), .A2(new_n448_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n451_), .A2(new_n452_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT85), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n449_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n487_), .B(KEYINPUT4), .C1(new_n488_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT98), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n481_), .A2(new_n486_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT4), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n455_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G225gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT97), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n494_), .A2(new_n495_), .A3(new_n498_), .A4(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n455_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n487_), .A3(new_n499_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n498_), .A2(new_n500_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n495_), .B1(new_n505_), .B2(new_n494_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n462_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n494_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n500_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT98), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n462_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n503_), .A4(new_n501_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n458_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n516_));
  AND4_X1   g315(.A1(new_n515_), .A2(new_n481_), .A3(new_n516_), .A4(new_n486_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n488_), .B2(new_n516_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G22gat), .B(G50gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n517_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n481_), .A2(new_n516_), .A3(new_n486_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT28), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n488_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n519_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT93), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G78gat), .B(G106gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT93), .B(new_n529_), .C1(new_n521_), .C2(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n533_));
  INV_X1    g332(.A(G204gat), .ZN(new_n534_));
  INV_X1    g333(.A(G197gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT90), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G197gat), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n534_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(G197gat), .A2(G204gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n533_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G218gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G211gat), .ZN(new_n543_));
  INV_X1    g342(.A(G211gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(G218gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n536_), .A2(new_n538_), .A3(new_n534_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT21), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(G197gat), .B2(G204gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n546_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n539_), .A2(new_n540_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n548_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n555_), .B(KEYINPUT92), .C1(new_n488_), .C2(new_n516_), .ZN(new_n556_));
  INV_X1    g355(.A(G233gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n488_), .A2(new_n516_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n541_), .A2(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n562_), .B(new_n560_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n520_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n523_), .A2(new_n524_), .A3(new_n519_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n532_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n532_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n531_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n566_), .A2(new_n567_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT94), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n579_), .A2(new_n574_), .A3(new_n528_), .A4(new_n530_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G226gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT19), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n404_), .A2(new_n405_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n427_), .A2(new_n408_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n394_), .A2(new_n419_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n423_), .A2(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT95), .B1(new_n588_), .B2(new_n564_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT25), .B(G183gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(G190gat), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n590_), .A2(new_n591_), .B1(new_n421_), .B2(new_n417_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n592_), .A2(new_n420_), .A3(new_n405_), .A4(new_n404_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n587_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n555_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n428_), .B2(new_n564_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n584_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G8gat), .B(G36gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT18), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G64gat), .B(G92gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n428_), .A2(new_n564_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n595_), .A2(new_n555_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n584_), .A2(KEYINPUT20), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n601_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT27), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n588_), .A2(new_n564_), .A3(KEYINPUT95), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n596_), .B1(new_n595_), .B2(new_n555_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n600_), .B(new_n584_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n595_), .B2(new_n555_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n583_), .B1(new_n607_), .B2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n605_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n611_), .A2(new_n612_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n608_), .A2(new_n609_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n607_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n395_), .A2(new_n398_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n419_), .A3(new_n409_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n423_), .A2(new_n427_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n564_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT20), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n589_), .B2(new_n597_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n605_), .B(new_n623_), .C1(new_n629_), .C2(new_n584_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT96), .ZN(new_n631_));
  INV_X1    g430(.A(new_n601_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n605_), .A4(new_n623_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n606_), .B1(new_n601_), .B2(new_n610_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n620_), .B1(new_n636_), .B2(new_n612_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n514_), .A2(new_n581_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n513_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n637_), .A2(new_n639_), .A3(new_n580_), .A4(new_n576_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n605_), .A2(KEYINPUT32), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n601_), .A2(new_n610_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n513_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT33), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n512_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n501_), .A2(new_n503_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(KEYINPUT33), .A3(new_n511_), .A4(new_n510_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n494_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n502_), .A2(new_n487_), .A3(new_n500_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n462_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT99), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n650_), .A2(new_n654_), .A3(new_n462_), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n647_), .A2(new_n649_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n645_), .B1(new_n657_), .B2(new_n636_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n581_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n640_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n638_), .B1(new_n660_), .B2(new_n458_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n316_), .A2(new_n369_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n367_), .A2(new_n368_), .A3(new_n309_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(G229gat), .A2(G233gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT78), .ZN(new_n666_));
  INV_X1    g465(.A(new_n309_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n368_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n365_), .B1(new_n357_), .B2(new_n363_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n663_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n664_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT78), .B(new_n664_), .C1(new_n670_), .C2(new_n663_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n665_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(G113gat), .B(G141gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT79), .ZN(new_n677_));
  XNOR2_X1  g476(.A(G169gat), .B(G197gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n665_), .B(new_n679_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(KEYINPUT80), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT80), .B1(new_n681_), .B2(new_n682_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n388_), .B1(new_n661_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n685_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n457_), .B1(new_n640_), .B2(new_n659_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT101), .B(new_n687_), .C1(new_n688_), .C2(new_n638_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n387_), .B1(new_n686_), .B2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n360_), .A3(new_n513_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT38), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n385_), .A2(new_n335_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n661_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n300_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n697_), .A2(KEYINPUT102), .A3(new_n685_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n300_), .B2(new_n687_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n383_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n698_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n696_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G1gat), .B1(new_n703_), .B2(new_n639_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n691_), .A2(new_n692_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n693_), .A2(new_n704_), .A3(new_n705_), .ZN(G1324gat));
  INV_X1    g505(.A(new_n637_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n690_), .A2(new_n361_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G8gat), .B1(new_n703_), .B2(new_n637_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT39), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT39), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n703_), .B2(new_n458_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n715_), .ZN(new_n717_));
  INV_X1    g516(.A(G15gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n690_), .A2(new_n718_), .A3(new_n457_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .ZN(G1326gat));
  OAI21_X1  g519(.A(G22gat), .B1(new_n703_), .B2(new_n581_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT42), .ZN(new_n722_));
  INV_X1    g521(.A(G22gat), .ZN(new_n723_));
  INV_X1    g522(.A(new_n581_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n690_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1327gat));
  NOR2_X1   g525(.A1(new_n383_), .A2(new_n694_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n300_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n686_), .B2(new_n689_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G29gat), .B1(new_n729_), .B2(new_n513_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n698_), .A2(new_n700_), .A3(new_n383_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n344_), .A2(new_n386_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n661_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n733_), .C1(new_n688_), .C2(new_n638_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n732_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT104), .B1(new_n738_), .B2(KEYINPUT44), .ZN(new_n739_));
  INV_X1    g538(.A(new_n737_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n514_), .A2(new_n637_), .A3(new_n581_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n576_), .A2(new_n639_), .A3(new_n580_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n742_), .A2(new_n637_), .B1(new_n658_), .B2(new_n581_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n743_), .B2(new_n457_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n736_), .B1(new_n744_), .B2(new_n733_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n731_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n739_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT44), .B(new_n731_), .C1(new_n740_), .C2(new_n745_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n738_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n750_), .A2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n513_), .A2(G29gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n730_), .B1(new_n756_), .B2(new_n757_), .ZN(G1328gat));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n750_), .A2(new_n755_), .A3(new_n707_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(G36gat), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n759_), .A2(new_n760_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n686_), .A2(new_n689_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n728_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n637_), .A2(G36gat), .ZN(new_n769_));
  AND4_X1   g568(.A1(new_n766_), .A2(new_n767_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n729_), .B2(new_n769_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n762_), .B1(new_n764_), .B2(new_n773_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n761_), .B(new_n772_), .C1(new_n763_), .C2(G36gat), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1329gat));
  NAND4_X1  g575(.A1(new_n750_), .A2(new_n755_), .A3(G43gat), .A4(new_n457_), .ZN(new_n777_));
  INV_X1    g576(.A(G43gat), .ZN(new_n778_));
  INV_X1    g577(.A(new_n729_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n458_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT47), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n777_), .A2(new_n783_), .A3(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1330gat));
  NAND3_X1  g584(.A1(new_n750_), .A2(new_n755_), .A3(new_n724_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(G50gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G50gat), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n581_), .A2(G50gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT108), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n788_), .A2(new_n789_), .B1(new_n779_), .B2(new_n791_), .ZN(G1331gat));
  NAND4_X1  g591(.A1(new_n696_), .A2(new_n685_), .A3(new_n697_), .A4(new_n383_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n793_), .A2(new_n238_), .A3(new_n639_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n661_), .A2(new_n687_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n733_), .A2(new_n300_), .A3(new_n701_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n639_), .B1(new_n797_), .B2(KEYINPUT109), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(KEYINPUT109), .B2(new_n797_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n794_), .B1(new_n799_), .B2(new_n238_), .ZN(G1332gat));
  OAI21_X1  g599(.A(G64gat), .B1(new_n793_), .B2(new_n637_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n797_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n236_), .A3(new_n707_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1333gat));
  OAI21_X1  g605(.A(G71gat), .B1(new_n793_), .B2(new_n458_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT49), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n457_), .A2(new_n246_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT111), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n797_), .B2(new_n810_), .ZN(G1334gat));
  OAI21_X1  g610(.A(G78gat), .B1(new_n793_), .B2(new_n581_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT50), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n804_), .A2(new_n244_), .A3(new_n724_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1335gat));
  NAND3_X1  g614(.A1(new_n795_), .A2(new_n697_), .A3(new_n727_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G85gat), .B1(new_n817_), .B2(new_n513_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n697_), .A2(new_n685_), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n383_), .B(new_n819_), .C1(new_n735_), .C2(new_n737_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT112), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n513_), .A2(new_n226_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(G1336gat));
  NAND3_X1  g622(.A1(new_n817_), .A2(new_n227_), .A3(new_n707_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n821_), .A2(new_n707_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n227_), .ZN(G1337gat));
  AOI21_X1  g625(.A(new_n213_), .B1(new_n820_), .B2(new_n457_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n457_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n817_), .B2(new_n828_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g629(.A1(new_n817_), .A2(new_n214_), .A3(new_n724_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n820_), .A2(new_n724_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(G106gat), .ZN(new_n834_));
  AOI211_X1 g633(.A(KEYINPUT52), .B(new_n214_), .C1(new_n820_), .C2(new_n724_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT53), .ZN(G1339gat));
  AND3_X1   g636(.A1(new_n344_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT54), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n838_), .A2(new_n685_), .A3(new_n300_), .A4(new_n840_), .ZN(new_n841_));
  XOR2_X1   g640(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n387_), .B2(new_n687_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n841_), .A2(new_n843_), .A3(KEYINPUT114), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT114), .B1(new_n841_), .B2(new_n843_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n295_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n283_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT55), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n283_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n281_), .A2(new_n282_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT12), .B1(new_n235_), .B2(new_n258_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n205_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT116), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n205_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n850_), .A2(new_n852_), .A3(new_n856_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n293_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(KEYINPUT56), .A3(new_n293_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n847_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n662_), .A2(new_n663_), .A3(new_n672_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n671_), .A2(new_n664_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n680_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n682_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n869_));
  OAI211_X1 g668(.A(KEYINPUT57), .B(new_n694_), .C1(new_n864_), .C2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n694_), .B1(new_n864_), .B2(new_n869_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n684_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n681_), .A2(KEYINPUT80), .A3(new_n682_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n289_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n859_), .A2(KEYINPUT56), .A3(new_n293_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n859_), .B2(new_n293_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n869_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n883_), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n694_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n289_), .A2(new_n868_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT58), .B(new_n885_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n733_), .A3(new_n889_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n872_), .A2(new_n875_), .A3(new_n884_), .A4(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n846_), .B1(new_n891_), .B2(new_n701_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n637_), .A2(new_n581_), .A3(new_n513_), .A4(new_n457_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n446_), .A3(new_n687_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n894_), .A2(KEYINPUT59), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(KEYINPUT59), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n685_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n895_), .B1(new_n898_), .B2(new_n446_), .ZN(G1340gat));
  OAI21_X1  g698(.A(new_n444_), .B1(new_n300_), .B2(KEYINPUT60), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n894_), .B(new_n900_), .C1(KEYINPUT60), .C2(new_n444_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n300_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n444_), .ZN(G1341gat));
  AOI21_X1  g702(.A(G127gat), .B1(new_n894_), .B2(new_n383_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n896_), .A2(new_n897_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n383_), .A2(G127gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT118), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n905_), .B2(new_n907_), .ZN(G1342gat));
  AOI21_X1  g707(.A(G134gat), .B1(new_n894_), .B2(new_n695_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n733_), .A2(G134gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT119), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n905_), .B2(new_n911_), .ZN(G1343gat));
  NAND2_X1  g711(.A1(new_n891_), .A2(new_n701_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n846_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NOR4_X1   g714(.A1(new_n707_), .A2(new_n581_), .A3(new_n639_), .A4(new_n457_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT120), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(KEYINPUT120), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G141gat), .B1(new_n921_), .B2(new_n685_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n463_), .B(new_n687_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1344gat));
  OAI21_X1  g723(.A(G148gat), .B1(new_n921_), .B2(new_n300_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n464_), .B(new_n697_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1345gat));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n921_), .B2(new_n701_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n928_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n383_), .B(new_n930_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1346gat));
  INV_X1    g731(.A(new_n920_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n734_), .B1(new_n933_), .B2(new_n918_), .ZN(new_n934_));
  INV_X1    g733(.A(G162gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n695_), .A2(new_n935_), .ZN(new_n936_));
  OAI22_X1  g735(.A1(new_n934_), .A2(new_n935_), .B1(new_n921_), .B2(new_n936_), .ZN(G1347gat));
  AND2_X1   g736(.A1(new_n687_), .A2(new_n396_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n707_), .A2(new_n514_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n940_), .A2(KEYINPUT121), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(KEYINPUT121), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n941_), .A2(new_n581_), .A3(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n939_), .B1(new_n915_), .B2(new_n944_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n892_), .A2(KEYINPUT123), .A3(new_n943_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n938_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n943_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n949_));
  AOI211_X1 g748(.A(new_n389_), .B(new_n948_), .C1(new_n949_), .C2(new_n687_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n948_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n915_), .A2(new_n687_), .A3(new_n944_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(G169gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n947_), .B1(new_n950_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(KEYINPUT124), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956_));
  OAI211_X1 g755(.A(new_n947_), .B(new_n956_), .C1(new_n950_), .C2(new_n953_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n955_), .A2(new_n957_), .ZN(G1348gat));
  OR2_X1    g757(.A1(new_n945_), .A2(new_n946_), .ZN(new_n959_));
  AOI21_X1  g758(.A(G176gat), .B1(new_n959_), .B2(new_n697_), .ZN(new_n960_));
  NOR4_X1   g759(.A1(new_n892_), .A2(new_n393_), .A3(new_n300_), .A4(new_n943_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962_));
  OR2_X1    g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n962_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n960_), .B1(new_n963_), .B2(new_n964_), .ZN(G1349gat));
  AOI21_X1  g764(.A(G183gat), .B1(new_n949_), .B2(new_n383_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n701_), .A2(new_n590_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n959_), .B2(new_n967_), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n959_), .A2(new_n591_), .A3(new_n695_), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n959_), .A2(new_n733_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n969_), .B1(new_n970_), .B2(new_n407_), .ZN(G1351gat));
  NAND3_X1  g770(.A1(new_n707_), .A2(new_n742_), .A3(new_n458_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n892_), .A2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(new_n687_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n697_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g776(.A1(new_n973_), .A2(new_n383_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n979_));
  AND2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n978_), .A2(new_n979_), .A3(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n978_), .B2(new_n979_), .ZN(G1354gat));
  XNOR2_X1  g781(.A(KEYINPUT126), .B(G218gat), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n973_), .A2(new_n733_), .A3(new_n983_), .ZN(new_n984_));
  NOR3_X1   g783(.A1(new_n892_), .A2(new_n694_), .A3(new_n972_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n984_), .B1(new_n985_), .B2(new_n983_), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n986_), .B(new_n987_), .ZN(G1355gat));
endmodule


