//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n202_));
  INV_X1    g001(.A(G57gat), .ZN(new_n203_));
  INV_X1    g002(.A(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G57gat), .A2(G64gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n202_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n202_), .A3(new_n206_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n208_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n210_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n207_), .A3(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G85gat), .B(G92gat), .Z(new_n230_));
  OAI211_X1 g029(.A(new_n226_), .B(new_n229_), .C1(new_n230_), .C2(new_n228_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n227_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n222_), .B(KEYINPUT6), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(KEYINPUT65), .A3(new_n236_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT8), .A3(new_n230_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n236_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n230_), .B1(new_n224_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT8), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n234_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n219_), .A2(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n219_), .A2(new_n251_), .A3(KEYINPUT67), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n234_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n214_), .A2(new_n218_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n252_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n251_), .A2(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n221_), .A2(new_n224_), .A3(new_n232_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n264_), .A2(new_n231_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT68), .B1(new_n265_), .B2(new_n246_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT12), .B(new_n219_), .C1(new_n263_), .C2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n260_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n252_), .B2(new_n271_), .ZN(new_n272_));
  AOI211_X1 g071(.A(KEYINPUT70), .B(new_n270_), .C1(new_n219_), .C2(new_n251_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n267_), .B(new_n268_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n261_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n279_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n261_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n282_), .A2(KEYINPUT71), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(new_n282_), .B2(KEYINPUT71), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n280_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(KEYINPUT71), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT72), .ZN(new_n288_));
  INV_X1    g087(.A(new_n280_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(KEYINPUT71), .A3(new_n283_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n286_), .A2(new_n291_), .A3(KEYINPUT13), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT13), .B1(new_n286_), .B2(new_n291_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT73), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G1gat), .B(G8gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G15gat), .ZN(new_n300_));
  INV_X1    g099(.A(G22gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G15gat), .A2(G22gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G1gat), .A2(G8gat), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n302_), .A2(new_n303_), .B1(KEYINPUT14), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n299_), .B(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G43gat), .B(G50gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(G29gat), .B(G36gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n296_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n299_), .A2(new_n305_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n299_), .A2(new_n305_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n311_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(KEYINPUT80), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G229gat), .A2(G233gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n311_), .B(KEYINPUT15), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n306_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n312_), .A2(new_n317_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n322_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G169gat), .B(G197gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n322_), .B(new_n329_), .C1(new_n319_), .C2(new_n323_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n295_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G204gat), .ZN(new_n333_));
  AND2_X1   g132(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G197gat), .A2(G204gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT21), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(G204gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT21), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(G197gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n338_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n341_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT91), .B(G197gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(G204gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT92), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT21), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n339_), .A2(new_n349_), .A3(new_n341_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n343_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n350_), .A2(new_n353_), .A3(KEYINPUT93), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT93), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n343_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n339_), .A2(new_n341_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n340_), .B1(new_n357_), .B2(KEYINPUT92), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n345_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G176gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT82), .B(new_n361_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n366_), .A2(new_n367_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT26), .B(G190gat), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT25), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(G183gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT81), .B1(new_n376_), .B2(KEYINPUT25), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n375_), .A2(new_n377_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n383_));
  AND3_X1   g182(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n368_), .ZN(new_n385_));
  OR2_X1    g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT24), .A3(new_n367_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n374_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n360_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT93), .B1(new_n350_), .B2(new_n353_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n356_), .A2(new_n358_), .A3(new_n355_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n344_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n379_), .A2(G183gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n375_), .A2(new_n377_), .A3(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n372_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n390_), .A2(KEYINPUT20), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(KEYINPUT98), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n390_), .A2(KEYINPUT20), .A3(new_n399_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n403_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  AOI211_X1 g208(.A(new_n344_), .B(new_n389_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT96), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n393_), .A2(new_n398_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT96), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(KEYINPUT20), .C1(new_n360_), .C2(new_n389_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n416_), .A2(KEYINPUT97), .A3(new_n407_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT97), .B1(new_n416_), .B2(new_n407_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n409_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420_));
  INV_X1    g219(.A(G92gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT18), .B(G64gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n426_), .B(new_n409_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n427_));
  INV_X1    g226(.A(G155gat), .ZN(new_n428_));
  INV_X1    g227(.A(G162gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT1), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(G155gat), .A3(G162gat), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n432_), .C1(G155gat), .C2(G162gat), .ZN(new_n433_));
  INV_X1    g232(.A(G141gat), .ZN(new_n434_));
  INV_X1    g233(.A(G148gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT3), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT3), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n442_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT2), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n441_), .A2(new_n443_), .A3(new_n445_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448_));
  XOR2_X1   g247(.A(G155gat), .B(G162gat), .Z(new_n449_));
  AND3_X1   g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n438_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT84), .B(G113gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G127gat), .B(G134gat), .ZN(new_n455_));
  INV_X1    g254(.A(G120gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n455_), .A2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n454_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n457_), .A3(new_n453_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n452_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT99), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n452_), .A2(new_n464_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n463_), .B(new_n438_), .C1(new_n451_), .C2(new_n450_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT4), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n472_), .B(KEYINPUT100), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT99), .A4(KEYINPUT4), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G29gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G85gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT0), .B(G57gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n468_), .A2(new_n469_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n473_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n476_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n471_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n474_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n480_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT33), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n485_), .A2(new_n489_), .A3(new_n480_), .A4(new_n486_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n484_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n425_), .A2(new_n427_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT101), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n486_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n481_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n487_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT102), .B1(new_n400_), .B2(new_n403_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n412_), .A2(new_n403_), .A3(new_n415_), .A4(new_n413_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT102), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n406_), .A2(new_n500_), .A3(new_n407_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n497_), .B(new_n504_), .C1(new_n419_), .C2(new_n503_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n425_), .A2(new_n491_), .A3(KEYINPUT101), .A4(new_n427_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n494_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G78gat), .B(G106gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G22gat), .B(G50gat), .Z(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n514_));
  INV_X1    g313(.A(new_n438_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n447_), .A2(new_n449_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT87), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n514_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G233gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n452_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n521_), .A2(new_n527_), .A3(new_n360_), .A4(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n519_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n531_), .B2(new_n393_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n519_), .A2(new_n520_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n513_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(new_n532_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n540_), .A2(new_n541_), .A3(new_n512_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT83), .B(G71gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT30), .B(G15gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n389_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n374_), .A2(new_n388_), .A3(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G227gat), .A2(G233gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(G99gat), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n547_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT85), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n464_), .A2(KEYINPUT31), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT31), .B1(new_n460_), .B2(new_n462_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n550_), .A2(new_n551_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n553_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n547_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n555_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n558_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n463_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT85), .B1(new_n571_), .B2(new_n561_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n558_), .B2(new_n567_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n545_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n507_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT27), .B1(new_n425_), .B2(new_n427_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n497_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n536_), .A2(new_n542_), .A3(new_n575_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n575_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n502_), .A2(new_n424_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n427_), .A2(KEYINPUT27), .A3(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n578_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n577_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n320_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n255_), .A2(new_n316_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n589_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n429_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT75), .B(G134gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n603_), .B(KEYINPUT36), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT37), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(KEYINPUT37), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n614_));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G183gat), .B(G211gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT78), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(G231gat), .A3(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(G231gat), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n619_), .B(new_n620_), .C1(new_n623_), .C2(new_n522_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n306_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n306_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n256_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n627_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n219_), .A3(new_n625_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT79), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n628_), .A2(new_n630_), .A3(KEYINPUT79), .A4(new_n631_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n612_), .A2(new_n613_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n332_), .A2(new_n587_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT103), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n332_), .A2(new_n639_), .A3(new_n587_), .A4(new_n636_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(G1gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n497_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n331_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n294_), .A2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT104), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT104), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n585_), .B1(new_n507_), .B2(new_n576_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n634_), .A2(new_n635_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n651_), .A2(new_n653_), .A3(new_n610_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n579_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n641_), .A2(KEYINPUT38), .A3(new_n642_), .A4(new_n497_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n656_), .A3(new_n657_), .ZN(G1324gat));
  INV_X1    g457(.A(G8gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n578_), .A2(new_n584_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n638_), .A2(new_n659_), .A3(new_n661_), .A4(new_n640_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  INV_X1    g462(.A(new_n655_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n661_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n665_), .B2(G8gat), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT39), .B(new_n659_), .C1(new_n664_), .C2(new_n661_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT40), .B(new_n662_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(new_n575_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G15gat), .B1(new_n655_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT41), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n641_), .A2(new_n300_), .A3(new_n575_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1326gat));
  NAND3_X1  g476(.A1(new_n641_), .A2(new_n301_), .A3(new_n545_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G22gat), .B1(new_n655_), .B2(new_n544_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT42), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n612_), .A2(new_n613_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n577_), .B2(new_n586_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n651_), .A2(KEYINPUT105), .A3(KEYINPUT43), .A4(new_n684_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n684_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(new_n587_), .B2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n687_), .A2(new_n688_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n650_), .A2(new_n653_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n682_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n587_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n651_), .B2(new_n684_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n685_), .A2(new_n683_), .A3(new_n686_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n652_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(new_n497_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G29gat), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n653_), .A2(new_n610_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n647_), .A2(new_n651_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n579_), .A2(G29gat), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT106), .Z(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n705_), .B2(new_n707_), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n693_), .A2(new_n661_), .A3(new_n700_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n660_), .A2(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n705_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n704_), .A2(new_n714_), .A3(new_n711_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n713_), .A2(KEYINPUT45), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT45), .B1(new_n713_), .B2(new_n715_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n710_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n710_), .A2(KEYINPUT46), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n693_), .A2(G43gat), .A3(new_n575_), .A4(new_n700_), .ZN(new_n724_));
  INV_X1    g523(.A(G43gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n705_), .B2(new_n673_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n693_), .A2(new_n545_), .A3(new_n700_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n693_), .A2(KEYINPUT108), .A3(new_n545_), .A4(new_n700_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(G50gat), .A3(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n544_), .A2(G50gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n705_), .B2(new_n734_), .ZN(G1331gat));
  INV_X1    g534(.A(new_n295_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n646_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT111), .B(G57gat), .Z(new_n738_));
  NAND4_X1  g537(.A1(new_n737_), .A2(new_n497_), .A3(new_n654_), .A4(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT112), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n651_), .A2(KEYINPUT109), .A3(new_n646_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT109), .B1(new_n651_), .B2(new_n646_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n294_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n636_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT110), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n497_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n740_), .B1(new_n747_), .B2(new_n203_), .ZN(G1332gat));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n204_), .A3(new_n661_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n737_), .A2(new_n654_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G64gat), .B1(new_n750_), .B2(new_n660_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT48), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n754_), .A3(new_n575_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G71gat), .B1(new_n750_), .B2(new_n673_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT49), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n746_), .A2(new_n759_), .A3(new_n545_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G78gat), .B1(new_n750_), .B2(new_n544_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT50), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1335gat));
  INV_X1    g562(.A(new_n703_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n741_), .A2(new_n295_), .A3(new_n764_), .A4(new_n742_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n765_), .A2(new_n579_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n744_), .A2(new_n331_), .A3(new_n653_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n698_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT114), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n698_), .A2(new_n771_), .A3(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n497_), .ZN(new_n774_));
  MUX2_X1   g573(.A(new_n766_), .B(new_n774_), .S(G85gat), .Z(G1336gat));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n421_), .B(new_n660_), .C1(new_n770_), .C2(new_n772_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n421_), .B1(new_n765_), .B2(new_n660_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT115), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n778_), .B(KEYINPUT115), .Z(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(G92gat), .A3(new_n661_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(KEYINPUT116), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n769_), .B2(new_n673_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n786_));
  OR3_X1    g585(.A1(new_n765_), .A2(new_n220_), .A3(new_n673_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  OR2_X1    g587(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(G1338gat));
  OR3_X1    g589(.A1(new_n765_), .A2(G106gat), .A3(new_n544_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n698_), .A2(new_n545_), .A3(new_n768_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G106gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n791_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  NAND2_X1  g599(.A1(new_n660_), .A2(new_n497_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n580_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n319_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n318_), .A2(new_n804_), .A3(new_n321_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n804_), .B2(new_n323_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n330_), .B1(new_n806_), .B2(new_n329_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n282_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n331_), .A2(new_n811_), .ZN(new_n812_));
  OAI221_X1 g611(.A(new_n267_), .B1(new_n257_), .B2(new_n253_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n260_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n272_), .A2(new_n273_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n815_), .A2(KEYINPUT55), .A3(new_n267_), .A4(new_n268_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n274_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n279_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n812_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n810_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n609_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(KEYINPUT57), .A3(new_n609_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n819_), .A2(new_n279_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n811_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n809_), .B(new_n282_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n836_), .A3(new_n689_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n827_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT119), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n826_), .A2(new_n840_), .A3(new_n837_), .A4(new_n827_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n653_), .A3(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n636_), .B(new_n331_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n803_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847_), .B2(new_n646_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n646_), .B2(KEYINPUT121), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n842_), .A2(new_n846_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n803_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(KEYINPUT59), .A3(new_n852_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n852_), .A2(KEYINPUT120), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(KEYINPUT120), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n838_), .A2(new_n653_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n854_), .B(new_n855_), .C1(new_n856_), .C2(new_n845_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n850_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n849_), .A2(KEYINPUT121), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n848_), .B1(new_n860_), .B2(new_n861_), .ZN(G1340gat));
  OR2_X1    g661(.A1(new_n456_), .A2(KEYINPUT60), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n847_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n456_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(KEYINPUT122), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT122), .B1(new_n864_), .B2(new_n865_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n736_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n456_), .B2(new_n868_), .ZN(G1341gat));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n847_), .A2(new_n870_), .A3(new_n652_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n653_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n870_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT123), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n871_), .B(new_n875_), .C1(new_n872_), .C2(new_n870_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n847_), .B2(new_n610_), .ZN(new_n878_));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n689_), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n851_), .A2(new_n581_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n801_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n646_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n295_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g686(.A1(new_n851_), .A2(new_n652_), .A3(new_n581_), .A4(new_n802_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n888_), .A2(KEYINPUT124), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(KEYINPUT124), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n889_), .A2(new_n890_), .A3(new_n892_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  AOI21_X1  g695(.A(G162gat), .B1(new_n883_), .B2(new_n610_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n684_), .A2(new_n429_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT125), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n883_), .B2(new_n899_), .ZN(G1347gat));
  NAND3_X1  g699(.A1(new_n661_), .A2(new_n579_), .A3(new_n575_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n838_), .A2(new_n653_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n545_), .B(new_n901_), .C1(new_n846_), .C2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n646_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(G169gat), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n904_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n362_), .A2(new_n363_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n907_), .B(new_n908_), .C1(new_n909_), .C2(new_n904_), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n903_), .B2(new_n744_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n851_), .A2(new_n544_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT126), .ZN(new_n913_));
  INV_X1    g712(.A(new_n901_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n851_), .A2(new_n915_), .A3(new_n544_), .ZN(new_n916_));
  AND4_X1   g715(.A1(new_n295_), .A2(new_n913_), .A3(new_n914_), .A4(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n911_), .B1(new_n917_), .B2(G176gat), .ZN(G1349gat));
  NAND4_X1  g717(.A1(new_n913_), .A2(new_n652_), .A3(new_n914_), .A4(new_n916_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n653_), .B1(new_n377_), .B2(new_n394_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n919_), .A2(new_n376_), .B1(new_n903_), .B2(new_n920_), .ZN(G1350gat));
  INV_X1    g720(.A(new_n903_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G190gat), .B1(new_n922_), .B2(new_n684_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n903_), .A2(new_n610_), .A3(new_n375_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n661_), .A2(new_n579_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n882_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n331_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT127), .B(G197gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n928_), .B2(new_n931_), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n882_), .A2(new_n926_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n295_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n933_), .B(new_n652_), .C1(new_n936_), .C2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n927_), .A2(new_n653_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n936_), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n933_), .B2(new_n610_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n933_), .A2(G218gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n689_), .ZN(G1355gat));
endmodule


