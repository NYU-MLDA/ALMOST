//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_;
  OR2_X1    g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  OAI22_X1  g003(.A1(new_n202_), .A2(KEYINPUT3), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT98), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n202_), .A2(KEYINPUT98), .A3(KEYINPUT3), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n205_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT99), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT96), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n214_), .A2(KEYINPUT94), .A3(KEYINPUT1), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n215_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT94), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT95), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n222_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT95), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n215_), .A4(new_n220_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n202_), .A2(new_n204_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT97), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT97), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n231_), .A3(new_n228_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n216_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  INV_X1    g035(.A(KEYINPUT103), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n237_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n233_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n227_), .A2(new_n231_), .A3(new_n228_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n231_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n236_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT103), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT4), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT104), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n246_), .A2(KEYINPUT4), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(new_n250_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT104), .B1(new_n259_), .B2(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n248_), .A2(new_n253_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G1gat), .B(G29gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G85gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT0), .B(G57gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT33), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT105), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n267_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT105), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT33), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n266_), .B1(new_n248_), .B2(new_n254_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n252_), .A2(new_n253_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n275_), .B1(new_n259_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G226gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT19), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT20), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G190gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT25), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G183gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT25), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OR3_X1    g092(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n287_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G169gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT85), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(G169gat), .B2(G176gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT24), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n295_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n285_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n290_), .A2(new_n291_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT100), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n290_), .A2(new_n306_), .A3(KEYINPUT100), .A4(new_n291_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT101), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(KEYINPUT86), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT86), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G169gat), .A3(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT22), .B(G169gat), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n297_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n311_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n312_), .B1(new_n311_), .B2(new_n318_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n304_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G211gat), .B(G218gat), .Z(new_n323_));
  INV_X1    g122(.A(KEYINPUT21), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n325_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n323_), .A3(KEYINPUT21), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n281_), .B1(new_n322_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n316_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n296_), .A2(KEYINPUT22), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT89), .ZN(new_n335_));
  AOI21_X1  g134(.A(G176gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n335_), .B2(new_n334_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n296_), .A2(KEYINPUT22), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT90), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n333_), .B(new_n307_), .C1(new_n337_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT24), .B1(new_n298_), .B2(new_n300_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n292_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n298_), .A2(new_n300_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n293_), .B(KEYINPUT88), .C1(new_n344_), .C2(KEYINPUT24), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n301_), .B2(new_n333_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT24), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n348_), .A2(new_n316_), .A3(KEYINPUT87), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n343_), .B(new_n345_), .C1(new_n347_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n285_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT82), .B1(new_n285_), .B2(KEYINPUT25), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n282_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT83), .B1(new_n285_), .B2(KEYINPUT25), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT83), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n283_), .A3(G183gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n351_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n353_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n285_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n355_), .A2(new_n357_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(KEYINPUT84), .A3(new_n363_), .A4(new_n282_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n340_), .B1(new_n350_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT102), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n330_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n366_), .B2(new_n330_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n332_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n321_), .A2(new_n330_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT20), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n366_), .A2(new_n330_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n279_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n370_), .A2(new_n374_), .A3(new_n379_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n271_), .A2(new_n274_), .A3(new_n277_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n330_), .B1(new_n233_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT28), .B1(new_n245_), .B2(KEYINPUT29), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT28), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n233_), .A2(new_n388_), .A3(new_n385_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(G78gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G106gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G22gat), .B(G50gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OR3_X1    g198(.A1(new_n390_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n269_), .A2(KEYINPUT106), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT106), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n272_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n266_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n250_), .B1(new_n249_), .B2(new_n256_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n259_), .A2(new_n255_), .A3(KEYINPUT104), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n262_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n404_), .A2(new_n406_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n321_), .B2(new_n330_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n331_), .B(new_n340_), .C1(new_n365_), .C2(new_n350_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n280_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n366_), .A2(new_n330_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT102), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n366_), .A2(new_n367_), .A3(new_n330_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n419_), .B2(new_n332_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n372_), .A2(new_n279_), .A3(new_n373_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n330_), .B1(new_n303_), .B2(new_n295_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n311_), .A2(new_n318_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n412_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n279_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n422_), .B1(new_n428_), .B2(new_n421_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n384_), .B(new_n403_), .C1(new_n411_), .C2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n410_), .A2(new_n407_), .ZN(new_n431_));
  AOI211_X1 g230(.A(KEYINPUT106), .B(new_n267_), .C1(new_n260_), .C2(new_n257_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n405_), .B1(new_n261_), .B2(new_n268_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n381_), .A2(new_n435_), .A3(new_n382_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT107), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n280_), .B1(new_n419_), .B2(new_n426_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n437_), .B(new_n380_), .C1(new_n438_), .C2(new_n423_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT107), .B1(new_n420_), .B2(new_n379_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n427_), .A2(new_n279_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n423_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n379_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n436_), .B1(new_n444_), .B2(KEYINPUT27), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n402_), .B1(new_n434_), .B2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G71gat), .B(G99gat), .Z(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G43gat), .ZN(new_n448_));
  AND2_X1   g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT91), .B(G15gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n366_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n366_), .A2(new_n453_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n458_), .A2(new_n454_), .A3(new_n451_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n450_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n236_), .B(KEYINPUT31), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n463_), .B2(KEYINPUT92), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n451_), .B1(new_n458_), .B2(new_n454_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n455_), .A2(new_n456_), .A3(new_n452_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n450_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n460_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n464_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n430_), .A2(new_n446_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT109), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT108), .B1(new_n445_), .B2(new_n402_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT108), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n382_), .A2(new_n437_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n379_), .B2(new_n428_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n435_), .B1(new_n480_), .B2(new_n439_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n478_), .B(new_n403_), .C1(new_n481_), .C2(new_n436_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n431_), .B(new_n473_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n476_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  AOI211_X1 g285(.A(KEYINPUT109), .B(new_n484_), .C1(new_n477_), .C2(new_n482_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n475_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT65), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT10), .B(G99gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT64), .B(G106gat), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G85gat), .A3(G92gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(G85gat), .B(G92gat), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT9), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n494_), .A2(new_n497_), .A3(new_n499_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT7), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n494_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n493_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n503_), .B1(new_n508_), .B2(new_n500_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n502_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G29gat), .B(G36gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT73), .B1(new_n511_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n511_), .A2(KEYINPUT73), .A3(new_n516_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n510_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n522_), .A2(new_n523_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT70), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n526_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT76), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT77), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT74), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n526_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n518_), .A2(KEYINPUT74), .A3(new_n524_), .A4(new_n525_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n528_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(KEYINPUT75), .A3(new_n531_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT75), .B1(new_n544_), .B2(new_n531_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n533_), .B(new_n540_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n532_), .B1(new_n549_), .B2(new_n545_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n537_), .B(KEYINPUT36), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT78), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n548_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n488_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G230gat), .ZN(new_n557_));
  INV_X1    g356(.A(G233gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n510_), .A2(KEYINPUT66), .A3(KEYINPUT12), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n563_));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n560_), .B(new_n568_), .C1(KEYINPUT12), .C2(new_n510_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n510_), .A2(KEYINPUT66), .A3(KEYINPUT12), .A4(new_n567_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n559_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n559_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n510_), .B2(new_n567_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n567_), .B2(new_n510_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G120gat), .B(G148gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n581_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n572_), .A2(new_n575_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(KEYINPUT13), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G15gat), .B(G22gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G1gat), .A2(G8gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT14), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G1gat), .B(G8gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n527_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n595_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n516_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n516_), .B(new_n597_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n602_), .B2(new_n599_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT81), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G113gat), .B(G141gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT80), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n607_), .B(new_n608_), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n605_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n589_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n597_), .B(new_n567_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(KEYINPUT66), .A2(KEYINPUT17), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT17), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n621_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n617_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n624_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n617_), .B2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n614_), .A2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n556_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n411_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n548_), .B(new_n636_), .C1(new_n550_), .C2(new_n553_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(new_n629_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT79), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n488_), .A2(new_n613_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n642_), .A2(G1gat), .A3(new_n411_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT110), .A3(new_n634_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT110), .B1(new_n643_), .B2(new_n634_), .ZN(new_n645_));
  OAI221_X1 g444(.A(new_n633_), .B1(new_n634_), .B2(new_n643_), .C1(new_n644_), .C2(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n445_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n642_), .A2(G8gat), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n631_), .A2(new_n445_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G8gat), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(KEYINPUT39), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(KEYINPUT39), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n653_), .B(new_n655_), .ZN(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n632_), .B2(new_n474_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT41), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n642_), .A2(G15gat), .A3(new_n474_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1326gat));
  OAI21_X1  g459(.A(G22gat), .B1(new_n632_), .B2(new_n403_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n403_), .A2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n642_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(new_n629_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n555_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n641_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G29gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n434_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT114), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n488_), .A2(new_n672_), .A3(new_n638_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT112), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT112), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n488_), .A2(new_n675_), .A3(new_n672_), .A4(new_n638_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n488_), .A2(new_n638_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n676_), .A3(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n614_), .A2(new_n665_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT113), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n679_), .A2(KEYINPUT113), .A3(new_n680_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n679_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(new_n434_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n671_), .B1(new_n689_), .B2(G29gat), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT114), .B(new_n669_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n670_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n445_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n686_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n641_), .A2(new_n694_), .A3(new_n445_), .A4(new_n666_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT115), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(KEYINPUT115), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n702_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT45), .A3(new_n700_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n693_), .B1(new_n697_), .B2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n703_), .A2(new_n705_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT44), .B1(new_n681_), .B2(new_n682_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n695_), .B1(new_n709_), .B2(new_n685_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n708_), .B(KEYINPUT46), .C1(new_n710_), .C2(new_n694_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1329gat));
  AOI21_X1  g511(.A(G43gat), .B1(new_n668_), .B2(new_n473_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n687_), .A2(G43gat), .A3(new_n473_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n686_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n668_), .B2(new_n402_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n687_), .A2(G50gat), .A3(new_n402_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n686_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(new_n589_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n611_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n556_), .A2(new_n665_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n411_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n488_), .A2(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n640_), .A2(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n411_), .A2(G57gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n726_), .B2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n723_), .B2(new_n647_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT48), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n647_), .A2(G64gat), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT116), .Z(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n726_), .B2(new_n732_), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n723_), .B2(new_n474_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT49), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n474_), .A2(G71gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n726_), .B2(new_n736_), .ZN(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n723_), .B2(new_n403_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT50), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n402_), .A2(new_n393_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n726_), .B2(new_n740_), .ZN(G1335gat));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n679_), .A2(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n721_), .A2(new_n611_), .A3(new_n665_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n674_), .A2(new_n678_), .A3(KEYINPUT117), .A4(new_n676_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n411_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n725_), .A2(new_n666_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n411_), .A2(G85gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(G1336gat));
  OAI21_X1  g549(.A(G92gat), .B1(new_n746_), .B2(new_n647_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n647_), .A2(G92gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n748_), .B2(new_n752_), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n746_), .B2(new_n474_), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n748_), .A2(new_n495_), .A3(new_n474_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT51), .ZN(G1338gat));
  AND2_X1   g556(.A1(new_n744_), .A2(new_n402_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n395_), .B1(new_n679_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n748_), .A2(new_n496_), .A3(new_n403_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NOR2_X1   g566(.A1(new_n589_), .A2(new_n611_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(new_n635_), .A3(new_n637_), .A4(new_n665_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n569_), .A2(new_n559_), .A3(new_n570_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n572_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n572_), .A2(KEYINPUT118), .A3(new_n773_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n571_), .B2(KEYINPUT55), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n774_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n583_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n584_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n599_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n596_), .A2(new_n598_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n602_), .B2(new_n781_), .ZN(new_n783_));
  MUX2_X1   g582(.A(new_n603_), .B(new_n783_), .S(new_n609_), .Z(new_n784_));
  NAND2_X1  g583(.A1(new_n775_), .A2(new_n777_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n774_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n581_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n780_), .A2(KEYINPUT58), .A3(new_n784_), .A4(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n779_), .A2(new_n789_), .A3(new_n584_), .A4(new_n784_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n637_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n533_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n552_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n636_), .B1(new_n796_), .B2(new_n548_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n790_), .B(new_n793_), .C1(new_n794_), .C2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n779_), .A2(new_n789_), .A3(new_n611_), .A4(new_n584_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n784_), .A2(new_n585_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n555_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n555_), .A2(new_n801_), .A3(KEYINPUT57), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n798_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n665_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n798_), .A2(new_n804_), .A3(KEYINPUT119), .A4(new_n805_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n771_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n483_), .A2(new_n434_), .A3(new_n473_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n611_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n810_), .B2(new_n811_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n811_), .A2(KEYINPUT59), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n806_), .A2(new_n629_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n771_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT120), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n612_), .A2(KEYINPUT121), .ZN(new_n820_));
  MUX2_X1   g619(.A(KEYINPUT121), .B(new_n820_), .S(G113gat), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n813_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  OAI21_X1  g621(.A(G120gat), .B1(new_n818_), .B2(new_n721_), .ZN(new_n823_));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n721_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n812_), .B(new_n825_), .C1(KEYINPUT60), .C2(new_n824_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n812_), .B2(new_n665_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n665_), .A2(G127gat), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT122), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n819_), .B2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n812_), .B2(new_n554_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n638_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT123), .B(G134gat), .Z(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n819_), .B2(new_n835_), .ZN(G1343gat));
  NAND2_X1  g635(.A1(new_n808_), .A2(new_n809_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n771_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n403_), .A2(new_n473_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n841_), .A2(new_n411_), .A3(new_n445_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n612_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT124), .B(G141gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1344gat));
  INV_X1    g645(.A(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n589_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g648(.A1(new_n843_), .A2(new_n629_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT61), .B(G155gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  OR3_X1    g651(.A1(new_n843_), .A2(G162gat), .A3(new_n555_), .ZN(new_n853_));
  OAI21_X1  g652(.A(G162gat), .B1(new_n843_), .B2(new_n833_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1347gat));
  NOR2_X1   g654(.A1(new_n816_), .A2(new_n771_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n484_), .A2(new_n647_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n403_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n296_), .B1(new_n859_), .B2(new_n611_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT62), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n611_), .A3(new_n317_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(KEYINPUT62), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(G1348gat));
  AOI21_X1  g663(.A(G176gat), .B1(new_n859_), .B2(new_n589_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n810_), .A2(new_n402_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n589_), .A2(G176gat), .A3(new_n857_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1349gat));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n665_), .A3(new_n857_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n629_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n869_), .A2(new_n285_), .B1(new_n859_), .B2(new_n870_), .ZN(G1350gat));
  NAND3_X1  g670(.A1(new_n859_), .A2(new_n282_), .A3(new_n554_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n856_), .A2(new_n833_), .A3(new_n858_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n305_), .ZN(G1351gat));
  NOR3_X1   g673(.A1(new_n841_), .A2(new_n434_), .A3(new_n647_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT125), .B1(new_n839_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  INV_X1    g676(.A(new_n875_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n810_), .A2(new_n877_), .A3(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(G197gat), .B(new_n611_), .C1(new_n876_), .C2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT126), .ZN(new_n881_));
  INV_X1    g680(.A(G197gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n876_), .A2(new_n879_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n612_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n839_), .A2(KEYINPUT125), .A3(new_n875_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n877_), .B1(new_n810_), .B2(new_n878_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n887_), .A2(new_n888_), .A3(G197gat), .A4(new_n611_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n881_), .A2(new_n884_), .A3(new_n889_), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n887_), .A2(new_n589_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g691(.A(new_n629_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT63), .B(G211gat), .Z(new_n894_));
  AOI21_X1  g693(.A(KEYINPUT127), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n665_), .B(new_n894_), .C1(new_n876_), .C2(new_n879_), .ZN(new_n896_));
  OR2_X1    g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n893_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n898_), .B2(KEYINPUT127), .ZN(G1354gat));
  OR3_X1    g698(.A1(new_n883_), .A2(G218gat), .A3(new_n555_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G218gat), .B1(new_n883_), .B2(new_n833_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1355gat));
endmodule


