//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(G113gat), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT3), .Z(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n215_), .B(KEYINPUT2), .Z(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT1), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n210_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n213_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n219_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n217_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n209_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G225gat), .A2(G233gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n225_), .A2(KEYINPUT95), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT95), .B1(new_n225_), .B2(new_n228_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n209_), .A2(new_n224_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n229_), .A2(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n227_), .B1(new_n233_), .B2(new_n226_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT0), .B(G57gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(G85gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(G1gat), .B(G29gat), .Z(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G197gat), .B(G204gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT21), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT90), .Z(new_n248_));
  OR3_X1    g047(.A1(new_n244_), .A2(KEYINPUT89), .A3(KEYINPUT21), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT89), .B1(new_n244_), .B2(KEYINPUT21), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n245_), .A3(new_n250_), .A4(new_n246_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT23), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(G183gat), .A3(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  MUX2_X1   g056(.A(new_n257_), .B(new_n256_), .S(KEYINPUT82), .Z(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT24), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  MUX2_X1   g060(.A(new_n260_), .B(KEYINPUT24), .S(new_n261_), .Z(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT26), .B(G190gat), .Z(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT25), .B(G183gat), .Z(new_n264_));
  OAI211_X1 g063(.A(new_n258_), .B(new_n262_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n257_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT81), .B(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n259_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n252_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT79), .B(G183gat), .Z(new_n273_));
  OAI21_X1  g072(.A(new_n258_), .B1(G190gat), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT22), .B1(new_n275_), .B2(KEYINPUT80), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(KEYINPUT22), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n267_), .B(new_n276_), .C1(new_n277_), .C2(KEYINPUT80), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(new_n278_), .A3(new_n259_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n273_), .B2(KEYINPUT25), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n257_), .B(new_n262_), .C1(new_n281_), .C2(new_n263_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n272_), .B(KEYINPUT20), .C1(new_n283_), .C2(new_n252_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G226gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT19), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n252_), .A2(new_n271_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n252_), .B2(new_n283_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n288_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G8gat), .B(G36gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT93), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT94), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n288_), .A2(new_n292_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n293_), .A2(new_n302_), .A3(new_n300_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n271_), .B(KEYINPUT98), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(new_n252_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n287_), .B1(new_n310_), .B2(new_n291_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n284_), .A2(new_n286_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n301_), .B(KEYINPUT27), .C1(new_n300_), .C2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT83), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT30), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n283_), .B(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G15gat), .B(G43gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n323_), .A2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n317_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n329_));
  XOR2_X1   g128(.A(new_n209_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n323_), .A2(new_n324_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT85), .A3(new_n325_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n317_), .B(new_n330_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G22gat), .B(G50gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n252_), .A2(KEYINPUT88), .A3(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G78gat), .B(G106gat), .Z(new_n346_));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n345_), .B(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n342_), .A2(new_n343_), .A3(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n343_), .A2(new_n349_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n334_), .A2(new_n335_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n243_), .B(new_n316_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n300_), .A2(KEYINPUT32), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n293_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n242_), .B(new_n357_), .C1(new_n313_), .C2(new_n356_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n305_), .A2(new_n307_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n234_), .A2(KEYINPUT33), .A3(new_n239_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n233_), .A2(new_n226_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n225_), .B(KEYINPUT97), .Z(new_n362_));
  OAI211_X1 g161(.A(new_n361_), .B(new_n238_), .C1(new_n226_), .C2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n241_), .A2(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n359_), .A2(new_n360_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n334_), .A2(new_n335_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n352_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n355_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G230gat), .A2(G233gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT65), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT65), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT6), .ZN(new_n375_));
  AND2_X1   g174(.A1(G99gat), .A2(G106gat), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT10), .B(G99gat), .Z(new_n380_));
  INV_X1    g179(.A(G106gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G85gat), .B(G92gat), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT9), .ZN(new_n384_));
  NAND2_X1  g183(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(KEYINPUT9), .ZN(new_n386_));
  NOR2_X1   g185(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(G92gat), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n379_), .A2(new_n382_), .A3(new_n384_), .A4(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT68), .B(G71gat), .ZN(new_n390_));
  INV_X1    g189(.A(G78gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G57gat), .B(G64gat), .Z(new_n393_));
  INV_X1    g192(.A(KEYINPUT11), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n394_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n390_), .B(G78gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT8), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT67), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n376_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n374_), .A2(KEYINPUT6), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n372_), .A2(KEYINPUT65), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(KEYINPUT67), .A3(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT7), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n404_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n402_), .B1(new_n413_), .B2(new_n383_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT7), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n415_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n408_), .A3(new_n417_), .A4(new_n409_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n402_), .A3(new_n383_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n389_), .B(new_n401_), .C1(new_n414_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n389_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n401_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n371_), .B(new_n423_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n425_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n421_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n371_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G120gat), .B(G148gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G204gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT5), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(G176gat), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n438_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n439_), .B(new_n440_), .C1(KEYINPUT70), .C2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G8gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(G15gat), .B(G22gat), .Z(new_n448_));
  OR2_X1    g247(.A1(KEYINPUT75), .A2(G1gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(KEYINPUT75), .A2(G1gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(G8gat), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT14), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(KEYINPUT76), .A3(KEYINPUT14), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n448_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G1gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI211_X1 g257(.A(G1gat), .B(new_n448_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n447_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n455_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT76), .B1(new_n451_), .B2(KEYINPUT14), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(G1gat), .B1(new_n463_), .B2(new_n448_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(new_n457_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(G8gat), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(G43gat), .ZN(new_n470_));
  INV_X1    g269(.A(G50gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n469_), .A2(G43gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(G43gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(G50gat), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT15), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(KEYINPUT15), .A3(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n468_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n472_), .A2(new_n475_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n467_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n481_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n460_), .A2(new_n466_), .A3(new_n482_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n482_), .B1(new_n460_), .B2(new_n466_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT78), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(new_n203_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n485_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n446_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G232gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT71), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT34), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n483_), .B(new_n389_), .C1(new_n414_), .C2(new_n420_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n389_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n413_), .A2(new_n383_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT8), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n510_), .B2(new_n419_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n478_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(new_n476_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n506_), .B(new_n507_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n504_), .A2(new_n505_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n479_), .A2(new_n424_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(KEYINPUT73), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT72), .B(G190gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G218gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G134gat), .B(G162gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT36), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n516_), .A2(new_n519_), .A3(KEYINPUT73), .A4(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n516_), .A2(new_n519_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT36), .A3(new_n524_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT74), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT37), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(KEYINPUT37), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(KEYINPUT37), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n529_), .A2(new_n535_), .A3(new_n531_), .A4(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT77), .Z(new_n540_));
  XOR2_X1   g339(.A(new_n401_), .B(new_n540_), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(new_n467_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT16), .B(G183gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G211gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n542_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(KEYINPUT17), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n538_), .A2(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n370_), .A2(new_n501_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n449_), .A2(new_n450_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n242_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT38), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT99), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n556_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n551_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n532_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT100), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT100), .ZN(new_n563_));
  AOI211_X1 g362(.A(new_n563_), .B(new_n532_), .C1(new_n355_), .C2(new_n369_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n501_), .B(new_n560_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(G1gat), .B1(new_n565_), .B2(new_n243_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n558_), .A2(new_n559_), .A3(new_n566_), .ZN(G1324gat));
  NAND3_X1  g366(.A1(new_n553_), .A2(new_n447_), .A3(new_n315_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT39), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n561_), .B(KEYINPUT100), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(new_n315_), .A3(new_n501_), .A4(new_n560_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(G8gat), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n569_), .B(G8gat), .C1(new_n565_), .C2(new_n316_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n568_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(KEYINPUT40), .B(new_n568_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1325gat));
  OAI21_X1  g378(.A(G15gat), .B1(new_n565_), .B2(new_n368_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT41), .Z(new_n581_));
  INV_X1    g380(.A(G15gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n368_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n553_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(G1326gat));
  OAI21_X1  g384(.A(G22gat), .B1(new_n565_), .B2(new_n352_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT42), .ZN(new_n587_));
  INV_X1    g386(.A(G22gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n352_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n553_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(G1327gat));
  NOR3_X1   g390(.A1(new_n446_), .A2(new_n500_), .A3(new_n560_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT43), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n370_), .B2(new_n538_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n538_), .ZN(new_n595_));
  AOI211_X1 g394(.A(KEYINPUT43), .B(new_n595_), .C1(new_n355_), .C2(new_n369_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT44), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT44), .B(new_n592_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n242_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(G29gat), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n532_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n592_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n243_), .A2(G29gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(G1328gat));
  NAND3_X1  g409(.A1(new_n599_), .A2(new_n315_), .A3(new_n600_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(G36gat), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n608_), .A2(G36gat), .A3(new_n316_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT45), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT46), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n614_), .A3(KEYINPUT46), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1329gat));
  NAND4_X1  g418(.A1(new_n599_), .A2(G43gat), .A3(new_n583_), .A4(new_n600_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(KEYINPUT102), .A2(G43gat), .ZN(new_n621_));
  OR2_X1    g420(.A1(KEYINPUT102), .A2(G43gat), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n621_), .B(new_n622_), .C1(new_n608_), .C2(new_n368_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT47), .ZN(G1330gat));
  AND3_X1   g424(.A1(new_n599_), .A2(new_n589_), .A3(new_n600_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n589_), .A2(new_n471_), .ZN(new_n627_));
  OAI22_X1  g426(.A1(new_n626_), .A2(new_n471_), .B1(new_n608_), .B2(new_n627_), .ZN(G1331gat));
  NAND2_X1  g427(.A1(new_n552_), .A2(new_n446_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n370_), .B(new_n500_), .C1(new_n629_), .C2(KEYINPUT103), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(KEYINPUT103), .B2(new_n629_), .ZN(new_n631_));
  AOI21_X1  g430(.A(G57gat), .B1(new_n631_), .B2(new_n242_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n446_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n499_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n570_), .A2(new_n560_), .A3(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n243_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n632_), .B1(new_n636_), .B2(G57gat), .ZN(G1332gat));
  NAND4_X1  g436(.A1(new_n570_), .A2(new_n315_), .A3(new_n560_), .A4(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G64gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT104), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n641_), .A3(G64gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT48), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G64gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n631_), .A2(new_n646_), .A3(new_n315_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n640_), .A2(KEYINPUT48), .A3(new_n642_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(G1333gat));
  INV_X1    g448(.A(G71gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n631_), .A2(new_n650_), .A3(new_n583_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n635_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n652_), .B2(new_n583_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT49), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n653_), .A2(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n651_), .B1(new_n656_), .B2(new_n657_), .ZN(G1334gat));
  NAND4_X1  g457(.A1(new_n570_), .A2(new_n589_), .A3(new_n560_), .A4(new_n634_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G78gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT105), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n662_), .A3(G78gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT50), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n631_), .A2(new_n391_), .A3(new_n589_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(KEYINPUT50), .A3(new_n663_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(G1335gat));
  NOR3_X1   g468(.A1(new_n633_), .A2(new_n499_), .A3(new_n560_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n607_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G85gat), .B1(new_n671_), .B2(new_n242_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT106), .Z(new_n673_));
  OR2_X1    g472(.A1(new_n594_), .A2(new_n596_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n670_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n387_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n243_), .B1(new_n677_), .B2(new_n385_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n673_), .B1(new_n676_), .B2(new_n678_), .ZN(G1336gat));
  AOI21_X1  g478(.A(G92gat), .B1(new_n671_), .B2(new_n315_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n315_), .A2(G92gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n681_), .ZN(G1337gat));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(KEYINPUT51), .ZN(new_n684_));
  OAI21_X1  g483(.A(G99gat), .B1(new_n675_), .B2(new_n368_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n671_), .A2(new_n583_), .A3(new_n380_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n683_), .A2(KEYINPUT51), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1338gat));
  NAND3_X1  g488(.A1(new_n671_), .A2(new_n381_), .A3(new_n589_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n589_), .B(new_n670_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT52), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(new_n692_), .A3(G106gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n691_), .B2(G106gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g495(.A1(new_n315_), .A2(new_n243_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n353_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n534_), .A2(new_n500_), .A3(new_n537_), .A4(new_n560_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n700_), .A2(new_n446_), .A3(KEYINPUT108), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT108), .B1(new_n700_), .B2(new_n446_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT54), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT109), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n701_), .A3(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n486_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT112), .B1(new_n714_), .B2(new_n495_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n481_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n496_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n480_), .A2(new_n486_), .A3(new_n484_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(new_n498_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n429_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n426_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n430_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OR2_X1    g526(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n727_), .A2(new_n371_), .A3(new_n423_), .A4(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n432_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n723_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n438_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT56), .B1(new_n732_), .B2(new_n438_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n721_), .B(new_n439_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT58), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n732_), .A2(new_n438_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT56), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n438_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n742_), .A2(KEYINPUT58), .A3(new_n439_), .A4(new_n721_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n743_), .A3(new_n538_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n732_), .A2(KEYINPUT111), .A3(KEYINPUT56), .A4(new_n438_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n747_), .A2(new_n499_), .A3(new_n439_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n749_), .A3(new_n741_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n748_), .A2(new_n750_), .B1(new_n441_), .B2(new_n721_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n745_), .B(new_n746_), .C1(new_n751_), .C2(new_n532_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(new_n750_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n721_), .A2(new_n441_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n532_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT113), .B1(new_n755_), .B2(KEYINPUT57), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT57), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n744_), .B(new_n752_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n551_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n699_), .B1(new_n713_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT114), .ZN(new_n761_));
  AOI21_X1  g560(.A(G113gat), .B1(new_n761_), .B2(new_n499_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT59), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n698_), .B(KEYINPUT115), .Z(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT116), .B(new_n744_), .C1(new_n755_), .C2(KEYINPUT57), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n755_), .A2(KEYINPUT57), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n746_), .B1(new_n751_), .B2(new_n532_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT116), .B1(new_n768_), .B2(new_n744_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n560_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n708_), .A2(new_n712_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n763_), .B(new_n764_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT117), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n773_), .B(new_n776_), .C1(new_n760_), .C2(new_n763_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n500_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n762_), .B1(new_n778_), .B2(G113gat), .ZN(G1340gat));
  OAI211_X1 g578(.A(new_n773_), .B(new_n446_), .C1(new_n760_), .C2(new_n763_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT118), .B(G120gat), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n633_), .B2(KEYINPUT60), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n783_), .A2(KEYINPUT60), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n759_), .A2(new_n712_), .A3(new_n708_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n786_), .A2(KEYINPUT114), .A3(new_n698_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n786_), .B2(new_n698_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n784_), .B(new_n785_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT119), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n782_), .A2(new_n789_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1341gat));
  AOI21_X1  g593(.A(G127gat), .B1(new_n761_), .B2(new_n560_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n775_), .A2(new_n777_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n560_), .A2(G127gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT120), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n796_), .B2(new_n798_), .ZN(G1342gat));
  AOI21_X1  g598(.A(G134gat), .B1(new_n761_), .B2(new_n532_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n595_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G134gat), .ZN(G1343gat));
  NAND3_X1  g601(.A1(new_n786_), .A2(new_n354_), .A3(new_n697_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n500_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n633_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g606(.A1(new_n803_), .A2(new_n551_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  NOR2_X1   g609(.A1(new_n803_), .A2(new_n606_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(G162gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n803_), .A2(new_n595_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(G162gat), .B2(new_n813_), .ZN(G1347gat));
  NOR3_X1   g613(.A1(new_n316_), .A2(new_n368_), .A3(new_n242_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n499_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT121), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n352_), .B(new_n817_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G169gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT62), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n815_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n589_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n268_), .A3(new_n499_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1348gat));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n446_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n589_), .B1(new_n713_), .B2(new_n759_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n815_), .A2(G176gat), .A3(new_n446_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n825_), .A2(new_n267_), .B1(new_n826_), .B2(new_n827_), .ZN(G1349gat));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n560_), .A3(new_n815_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n273_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n560_), .A2(new_n264_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n829_), .A2(new_n830_), .B1(new_n822_), .B2(new_n831_), .ZN(G1350gat));
  NAND2_X1  g631(.A1(new_n822_), .A2(new_n538_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G190gat), .ZN(new_n834_));
  INV_X1    g633(.A(new_n263_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n822_), .A2(new_n835_), .A3(new_n532_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1351gat));
  NAND3_X1  g636(.A1(new_n354_), .A2(KEYINPUT122), .A3(new_n243_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT122), .B1(new_n354_), .B2(new_n243_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n316_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n786_), .A2(new_n838_), .A3(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n500_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(G197gat), .Z(G1352gat));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G204gat), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n841_), .A2(new_n633_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(G204gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n846_), .B2(new_n845_), .ZN(G1353gat));
  NAND4_X1  g648(.A1(new_n786_), .A2(new_n560_), .A3(new_n838_), .A4(new_n840_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT63), .B(G211gat), .Z(new_n851_));
  OR2_X1    g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n850_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1354gat));
  XNOR2_X1  g656(.A(KEYINPUT125), .B(G218gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n841_), .B2(new_n606_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n595_), .A2(new_n858_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n841_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1355gat));
endmodule


