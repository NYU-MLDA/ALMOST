//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_c1355" written by ABC on Sun Mar 26 01:26:03 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n508_, new_n509_, new_n510_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n556_, new_n557_, new_n558_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n671_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_;
  INV_X1    g000(.A(G183gat), .ZN(new_n138_));
  INV_X1    g001(.A(G190gat), .ZN(new_n139_));
  NAND2_X1  g002(.A1(new_n138_), .A2(new_n139_), .ZN(new_n140_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n141_));
  AOI21_X1  g004(.A(new_n141_), .B1(G183gat), .B2(G190gat), .ZN(new_n142_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n143_));
  NOR2_X1   g006(.A1(new_n143_), .A2(KEYINPUT23), .ZN(new_n144_));
  OAI21_X1  g007(.A(new_n140_), .B1(new_n142_), .B2(new_n144_), .ZN(new_n145_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n146_));
  XNOR2_X1  g009(.A(KEYINPUT22), .B(G169gat), .ZN(new_n147_));
  INV_X1    g010(.A(G176gat), .ZN(new_n148_));
  NAND2_X1  g011(.A1(new_n147_), .A2(new_n148_), .ZN(new_n149_));
  NAND3_X1  g012(.A1(new_n145_), .A2(new_n146_), .A3(new_n149_), .ZN(new_n150_));
  NAND2_X1  g013(.A1(new_n143_), .A2(KEYINPUT23), .ZN(new_n151_));
  NAND3_X1  g014(.A1(new_n141_), .A2(G183gat), .A3(G190gat), .ZN(new_n152_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n153_));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n154_));
  AOI22_X1  g017(.A1(new_n151_), .A2(new_n152_), .B1(new_n153_), .B2(new_n154_), .ZN(new_n155_));
  NAND2_X1  g018(.A1(new_n138_), .A2(KEYINPUT25), .ZN(new_n156_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n157_));
  NAND2_X1  g020(.A1(new_n157_), .A2(G183gat), .ZN(new_n158_));
  NAND2_X1  g021(.A1(new_n139_), .A2(KEYINPUT26), .ZN(new_n159_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n160_));
  NAND2_X1  g023(.A1(new_n160_), .A2(G190gat), .ZN(new_n161_));
  NAND4_X1  g024(.A1(new_n156_), .A2(new_n158_), .A3(new_n159_), .A4(new_n161_), .ZN(new_n162_));
  INV_X1    g025(.A(new_n154_), .ZN(new_n163_));
  NAND3_X1  g026(.A1(new_n163_), .A2(KEYINPUT24), .A3(new_n146_), .ZN(new_n164_));
  NAND3_X1  g027(.A1(new_n155_), .A2(new_n162_), .A3(new_n164_), .ZN(new_n165_));
  NAND2_X1  g028(.A1(new_n150_), .A2(new_n165_), .ZN(new_n166_));
  INV_X1    g029(.A(G134gat), .ZN(new_n167_));
  NAND2_X1  g030(.A1(new_n167_), .A2(G127gat), .ZN(new_n168_));
  INV_X1    g031(.A(G127gat), .ZN(new_n169_));
  NAND2_X1  g032(.A1(new_n169_), .A2(G134gat), .ZN(new_n170_));
  NAND2_X1  g033(.A1(new_n168_), .A2(new_n170_), .ZN(new_n171_));
  INV_X1    g034(.A(G120gat), .ZN(new_n172_));
  NAND2_X1  g035(.A1(new_n172_), .A2(G113gat), .ZN(new_n173_));
  INV_X1    g036(.A(G113gat), .ZN(new_n174_));
  NAND2_X1  g037(.A1(new_n174_), .A2(G120gat), .ZN(new_n175_));
  NAND2_X1  g038(.A1(new_n173_), .A2(new_n175_), .ZN(new_n176_));
  NAND2_X1  g039(.A1(new_n171_), .A2(new_n176_), .ZN(new_n177_));
  NAND4_X1  g040(.A1(new_n168_), .A2(new_n170_), .A3(new_n173_), .A4(new_n175_), .ZN(new_n178_));
  NAND2_X1  g041(.A1(new_n177_), .A2(new_n178_), .ZN(new_n179_));
  INV_X1    g042(.A(new_n179_), .ZN(new_n180_));
  XNOR2_X1  g043(.A(new_n166_), .B(new_n180_), .ZN(new_n181_));
  INV_X1    g044(.A(G71gat), .ZN(new_n182_));
  INV_X1    g045(.A(G99gat), .ZN(new_n183_));
  NAND2_X1  g046(.A1(new_n182_), .A2(new_n183_), .ZN(new_n184_));
  NAND2_X1  g047(.A1(G71gat), .A2(G99gat), .ZN(new_n185_));
  NAND2_X1  g048(.A1(new_n184_), .A2(new_n185_), .ZN(new_n186_));
  INV_X1    g049(.A(KEYINPUT31), .ZN(new_n187_));
  NAND2_X1  g050(.A1(new_n186_), .A2(new_n187_), .ZN(new_n188_));
  NAND3_X1  g051(.A1(new_n184_), .A2(KEYINPUT31), .A3(new_n185_), .ZN(new_n189_));
  NAND2_X1  g052(.A1(new_n188_), .A2(new_n189_), .ZN(new_n190_));
  NAND2_X1  g053(.A1(new_n190_), .A2(KEYINPUT30), .ZN(new_n191_));
  INV_X1    g054(.A(KEYINPUT30), .ZN(new_n192_));
  NAND3_X1  g055(.A1(new_n188_), .A2(new_n192_), .A3(new_n189_), .ZN(new_n193_));
  NAND4_X1  g056(.A1(new_n191_), .A2(G227gat), .A3(G233gat), .A4(new_n193_), .ZN(new_n194_));
  NAND2_X1  g057(.A1(G227gat), .A2(G233gat), .ZN(new_n195_));
  AND3_X1   g058(.A1(new_n188_), .A2(new_n192_), .A3(new_n189_), .ZN(new_n196_));
  AOI21_X1  g059(.A(new_n192_), .B1(new_n188_), .B2(new_n189_), .ZN(new_n197_));
  OAI21_X1  g060(.A(new_n195_), .B1(new_n196_), .B2(new_n197_), .ZN(new_n198_));
  XNOR2_X1  g061(.A(G15gat), .B(G43gat), .ZN(new_n199_));
  INV_X1    g062(.A(new_n199_), .ZN(new_n200_));
  AND3_X1   g063(.A1(new_n194_), .A2(new_n198_), .A3(new_n200_), .ZN(new_n201_));
  AOI21_X1  g064(.A(new_n200_), .B1(new_n194_), .B2(new_n198_), .ZN(new_n202_));
  OAI21_X1  g065(.A(new_n181_), .B1(new_n201_), .B2(new_n202_), .ZN(new_n203_));
  NAND2_X1  g066(.A1(new_n194_), .A2(new_n198_), .ZN(new_n204_));
  NAND2_X1  g067(.A1(new_n204_), .A2(new_n199_), .ZN(new_n205_));
  XNOR2_X1  g068(.A(new_n166_), .B(new_n179_), .ZN(new_n206_));
  NAND3_X1  g069(.A1(new_n194_), .A2(new_n198_), .A3(new_n200_), .ZN(new_n207_));
  NAND3_X1  g070(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AND2_X1   g071(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g072(.A(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n211_));
  INV_X1    g074(.A(KEYINPUT21), .ZN(new_n212_));
  NAND2_X1  g075(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g076(.A(G197gat), .ZN(new_n214_));
  NOR2_X1   g077(.A1(new_n214_), .A2(G204gat), .ZN(new_n215_));
  INV_X1    g078(.A(G204gat), .ZN(new_n216_));
  NOR2_X1   g079(.A1(new_n216_), .A2(G197gat), .ZN(new_n217_));
  OAI21_X1  g080(.A(KEYINPUT21), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n219_));
  NAND3_X1  g082(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n221_));
  OAI211_X1 g084(.A(new_n221_), .B(KEYINPUT21), .C1(new_n215_), .C2(new_n217_), .ZN(new_n222_));
  NAND2_X1  g085(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g086(.A(G78gat), .B(G106gat), .ZN(new_n224_));
  INV_X1    g087(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n226_));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n227_));
  INV_X1    g090(.A(G141gat), .ZN(new_n228_));
  INV_X1    g091(.A(G148gat), .ZN(new_n229_));
  NAND3_X1  g092(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n232_));
  NAND2_X1  g095(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g096(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  NAND3_X1  g097(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  NAND4_X1  g098(.A1(new_n230_), .A2(new_n233_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  OR2_X1    g099(.A1(G155gat), .A2(G162gat), .ZN(new_n237_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  AND2_X1   g101(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g102(.A1(new_n238_), .A2(KEYINPUT1), .ZN(new_n240_));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n241_));
  NAND3_X1  g104(.A1(new_n241_), .A2(G155gat), .A3(G162gat), .ZN(new_n242_));
  NAND3_X1  g105(.A1(new_n240_), .A2(new_n242_), .A3(new_n237_), .ZN(new_n243_));
  XOR2_X1   g106(.A(G141gat), .B(G148gat), .Z(new_n244_));
  AOI22_X1  g107(.A1(new_n236_), .A2(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g108(.A(new_n223_), .B(new_n225_), .C1(new_n226_), .C2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g109(.A(G22gat), .B(G50gat), .ZN(new_n247_));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n248_));
  XNOR2_X1  g111(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g112(.A(G228gat), .ZN(new_n250_));
  INV_X1    g113(.A(G233gat), .ZN(new_n251_));
  OAI21_X1  g114(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g115(.A(new_n247_), .B(KEYINPUT28), .ZN(new_n253_));
  NOR2_X1   g116(.A1(new_n250_), .A2(new_n251_), .ZN(new_n254_));
  NAND2_X1  g117(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g118(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g119(.A1(new_n236_), .A2(new_n239_), .ZN(new_n257_));
  NAND2_X1  g120(.A1(new_n243_), .A2(new_n244_), .ZN(new_n258_));
  NAND2_X1  g121(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g122(.A1(new_n259_), .A2(KEYINPUT29), .ZN(new_n260_));
  NAND2_X1  g123(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g124(.A(new_n223_), .B1(new_n226_), .B2(new_n245_), .ZN(new_n262_));
  NAND2_X1  g125(.A1(new_n262_), .A2(new_n224_), .ZN(new_n263_));
  OAI211_X1 g126(.A(new_n252_), .B(new_n255_), .C1(KEYINPUT29), .C2(new_n259_), .ZN(new_n264_));
  AND4_X1   g127(.A1(new_n246_), .A2(new_n261_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  AOI22_X1  g128(.A1(new_n261_), .A2(new_n264_), .B1(new_n263_), .B2(new_n246_), .ZN(new_n266_));
  NOR2_X1   g129(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g130(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g131(.A1(new_n166_), .A2(new_n223_), .ZN(new_n269_));
  NAND4_X1  g132(.A1(new_n150_), .A2(new_n220_), .A3(new_n165_), .A4(new_n222_), .ZN(new_n270_));
  NAND3_X1  g133(.A1(new_n269_), .A2(KEYINPUT20), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XOR2_X1   g135(.A(new_n272_), .B(KEYINPUT19), .Z(new_n273_));
  INV_X1    g136(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g137(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g138(.A1(new_n269_), .A2(KEYINPUT20), .A3(new_n273_), .A4(new_n270_), .ZN(new_n276_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n277_));
  XNOR2_X1  g140(.A(new_n277_), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g141(.A(KEYINPUT18), .B(G64gat), .ZN(new_n279_));
  XOR2_X1   g142(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  AND3_X1   g143(.A1(new_n275_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g144(.A(new_n280_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n282_));
  NOR2_X1   g145(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n285_));
  NAND2_X1  g148(.A1(new_n259_), .A2(new_n180_), .ZN(new_n286_));
  NAND2_X1  g149(.A1(new_n245_), .A2(new_n179_), .ZN(new_n287_));
  AOI21_X1  g150(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g151(.A1(new_n245_), .A2(new_n179_), .ZN(new_n289_));
  NOR2_X1   g152(.A1(new_n289_), .A2(KEYINPUT4), .ZN(new_n290_));
  OAI21_X1  g153(.A(new_n284_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n292_));
  XNOR2_X1  g155(.A(new_n292_), .B(G85gat), .ZN(new_n293_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n294_));
  XOR2_X1   g157(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  INV_X1    g158(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g159(.A(new_n284_), .ZN(new_n297_));
  NAND3_X1  g160(.A1(new_n286_), .A2(new_n297_), .A3(new_n287_), .ZN(new_n298_));
  NAND3_X1  g161(.A1(new_n291_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g162(.A(new_n297_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n300_));
  NAND3_X1  g163(.A1(new_n286_), .A2(new_n284_), .A3(new_n287_), .ZN(new_n301_));
  NAND3_X1  g164(.A1(new_n300_), .A2(new_n301_), .A3(new_n295_), .ZN(new_n302_));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n303_));
  NAND2_X1  g166(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g167(.A1(new_n300_), .A2(KEYINPUT33), .A3(new_n301_), .A4(new_n295_), .ZN(new_n305_));
  NAND4_X1  g168(.A1(new_n283_), .A2(new_n299_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g169(.A1(new_n280_), .A2(KEYINPUT32), .ZN(new_n307_));
  NAND3_X1  g170(.A1(new_n275_), .A2(new_n307_), .A3(new_n276_), .ZN(new_n308_));
  NAND2_X1  g171(.A1(new_n275_), .A2(new_n276_), .ZN(new_n309_));
  INV_X1    g172(.A(new_n307_), .ZN(new_n310_));
  NAND2_X1  g173(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AND3_X1   g174(.A1(new_n179_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n312_));
  OAI21_X1  g175(.A(KEYINPUT4), .B1(new_n312_), .B2(new_n289_), .ZN(new_n313_));
  NAND2_X1  g176(.A1(new_n286_), .A2(new_n285_), .ZN(new_n314_));
  AOI21_X1  g177(.A(new_n284_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g178(.A(new_n301_), .ZN(new_n316_));
  NOR3_X1   g179(.A1(new_n315_), .A2(new_n316_), .A3(new_n296_), .ZN(new_n317_));
  AOI21_X1  g180(.A(new_n295_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n318_));
  OAI211_X1 g181(.A(new_n308_), .B(new_n311_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g182(.A(new_n268_), .B1(new_n306_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g183(.A(new_n296_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n321_));
  NAND2_X1  g184(.A1(new_n321_), .A2(new_n302_), .ZN(new_n322_));
  OAI21_X1  g185(.A(KEYINPUT27), .B1(new_n281_), .B2(new_n282_), .ZN(new_n323_));
  INV_X1    g186(.A(new_n280_), .ZN(new_n324_));
  NAND2_X1  g187(.A1(new_n309_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n326_));
  NAND3_X1  g189(.A1(new_n275_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n327_));
  NAND3_X1  g190(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AOI211_X1 g191(.A(new_n267_), .B(new_n322_), .C1(new_n323_), .C2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g192(.A(new_n210_), .B1(new_n320_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g193(.A1(new_n209_), .A2(new_n321_), .A3(new_n302_), .ZN(new_n331_));
  INV_X1    g194(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g195(.A(new_n328_), .ZN(new_n333_));
  INV_X1    g196(.A(new_n323_), .ZN(new_n334_));
  OAI211_X1 g197(.A(new_n332_), .B(new_n267_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g198(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g199(.A1(G230gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g200(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g201(.A(KEYINPUT9), .ZN(new_n339_));
  INV_X1    g202(.A(G85gat), .ZN(new_n340_));
  INV_X1    g203(.A(G92gat), .ZN(new_n341_));
  OAI21_X1  g204(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g205(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n343_));
  OAI211_X1 g206(.A(new_n342_), .B(new_n343_), .C1(G85gat), .C2(G92gat), .ZN(new_n344_));
  NAND2_X1  g207(.A1(G99gat), .A2(G106gat), .ZN(new_n345_));
  NAND2_X1  g208(.A1(new_n345_), .A2(KEYINPUT6), .ZN(new_n346_));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n347_));
  NAND3_X1  g210(.A1(new_n347_), .A2(G99gat), .A3(G106gat), .ZN(new_n348_));
  NAND2_X1  g211(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  OR2_X1    g212(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n350_));
  INV_X1    g213(.A(G106gat), .ZN(new_n351_));
  NAND2_X1  g214(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n352_));
  NAND3_X1  g215(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AND3_X1   g216(.A1(new_n344_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g217(.A(G85gat), .B(G92gat), .ZN(new_n355_));
  INV_X1    g218(.A(new_n355_), .ZN(new_n356_));
  AND2_X1   g219(.A1(new_n346_), .A2(new_n348_), .ZN(new_n357_));
  INV_X1    g220(.A(KEYINPUT7), .ZN(new_n358_));
  NAND3_X1  g221(.A1(new_n358_), .A2(new_n183_), .A3(new_n351_), .ZN(new_n359_));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n360_));
  NAND2_X1  g223(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g224(.A(new_n356_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g225(.A1(new_n362_), .A2(KEYINPUT8), .ZN(new_n363_));
  NAND3_X1  g226(.A1(new_n349_), .A2(new_n360_), .A3(new_n359_), .ZN(new_n364_));
  INV_X1    g227(.A(KEYINPUT8), .ZN(new_n365_));
  NAND3_X1  g228(.A1(new_n364_), .A2(new_n365_), .A3(new_n356_), .ZN(new_n366_));
  AOI21_X1  g229(.A(new_n354_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g230(.A(G71gat), .B(G78gat), .Z(new_n368_));
  XNOR2_X1  g231(.A(G57gat), .B(G64gat), .ZN(new_n369_));
  OAI21_X1  g232(.A(new_n368_), .B1(KEYINPUT11), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g233(.A1(new_n369_), .A2(KEYINPUT11), .ZN(new_n371_));
  INV_X1    g234(.A(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g235(.A(new_n370_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g236(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g237(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g238(.A1(new_n367_), .A2(new_n373_), .ZN(new_n376_));
  OAI21_X1  g239(.A(new_n338_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n378_));
  OAI21_X1  g241(.A(new_n378_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n379_));
  AOI21_X1  g242(.A(new_n338_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n380_));
  NAND3_X1  g243(.A1(new_n344_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n381_));
  INV_X1    g244(.A(new_n360_), .ZN(new_n382_));
  NOR3_X1   g245(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n383_));
  NOR2_X1   g246(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI211_X1 g247(.A(KEYINPUT8), .B(new_n355_), .C1(new_n384_), .C2(new_n349_), .ZN(new_n385_));
  AOI21_X1  g248(.A(new_n365_), .B1(new_n364_), .B2(new_n356_), .ZN(new_n386_));
  OAI21_X1  g249(.A(new_n381_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g250(.A(new_n370_), .B(new_n371_), .ZN(new_n388_));
  NAND3_X1  g251(.A1(new_n387_), .A2(KEYINPUT12), .A3(new_n388_), .ZN(new_n389_));
  NAND3_X1  g252(.A1(new_n379_), .A2(new_n380_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g253(.A1(new_n377_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g254(.A(G120gat), .B(G148gat), .ZN(new_n392_));
  XNOR2_X1  g255(.A(new_n392_), .B(G204gat), .ZN(new_n393_));
  XNOR2_X1  g256(.A(KEYINPUT5), .B(G176gat), .ZN(new_n394_));
  XNOR2_X1  g257(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g258(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g259(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g260(.A1(new_n377_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n398_));
  NAND2_X1  g261(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g262(.A(KEYINPUT13), .ZN(new_n400_));
  NAND2_X1  g263(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g264(.A1(new_n397_), .A2(KEYINPUT13), .A3(new_n398_), .ZN(new_n402_));
  NAND2_X1  g265(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g266(.A(G29gat), .B(G36gat), .Z(new_n404_));
  XOR2_X1   g267(.A(G43gat), .B(G50gat), .Z(new_n405_));
  NAND2_X1  g268(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g269(.A(G29gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n408_));
  NAND2_X1  g271(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g272(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g273(.A(KEYINPUT15), .ZN(new_n411_));
  NAND2_X1  g274(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g275(.A1(new_n406_), .A2(KEYINPUT15), .A3(new_n409_), .ZN(new_n413_));
  NAND2_X1  g276(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n415_));
  INV_X1    g278(.A(G1gat), .ZN(new_n416_));
  INV_X1    g279(.A(G8gat), .ZN(new_n417_));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g281(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g282(.A(G1gat), .B(G8gat), .Z(new_n420_));
  XNOR2_X1  g283(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  OR2_X1    g284(.A1(new_n414_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n423_));
  NAND2_X1  g286(.A1(new_n421_), .A2(new_n410_), .ZN(new_n424_));
  NAND3_X1  g287(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g288(.A(new_n421_), .B(new_n410_), .ZN(new_n426_));
  NAND3_X1  g289(.A1(new_n426_), .A2(G229gat), .A3(G233gat), .ZN(new_n427_));
  NAND2_X1  g290(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n429_));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n430_));
  XOR2_X1   g293(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  INV_X1    g294(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g295(.A1(new_n428_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g296(.A1(new_n425_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n434_));
  AND2_X1   g297(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g298(.A1(new_n403_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g299(.A1(new_n336_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g300(.A(new_n437_), .ZN(new_n438_));
  OAI211_X1 g301(.A(new_n381_), .B(new_n410_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n439_));
  OAI21_X1  g302(.A(new_n439_), .B1(new_n367_), .B2(new_n414_), .ZN(new_n440_));
  NAND2_X1  g303(.A1(G232gat), .A2(G233gat), .ZN(new_n441_));
  XOR2_X1   g304(.A(new_n441_), .B(KEYINPUT34), .Z(new_n442_));
  INV_X1    g305(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g306(.A1(new_n440_), .A2(KEYINPUT35), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g307(.A1(new_n387_), .A2(new_n413_), .A3(new_n412_), .ZN(new_n445_));
  NAND2_X1  g308(.A1(new_n443_), .A2(KEYINPUT35), .ZN(new_n446_));
  OR2_X1    g309(.A1(new_n443_), .A2(KEYINPUT35), .ZN(new_n447_));
  NAND4_X1  g310(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(new_n439_), .ZN(new_n448_));
  AND3_X1   g311(.A1(new_n444_), .A2(new_n448_), .A3(KEYINPUT36), .ZN(new_n449_));
  AOI21_X1  g312(.A(KEYINPUT36), .B1(new_n444_), .B2(new_n448_), .ZN(new_n450_));
  XNOR2_X1  g313(.A(G134gat), .B(G162gat), .ZN(new_n451_));
  XNOR2_X1  g314(.A(G190gat), .B(G218gat), .ZN(new_n452_));
  XNOR2_X1  g315(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  NOR3_X1   g316(.A1(new_n449_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g317(.A1(new_n450_), .A2(new_n453_), .ZN(new_n455_));
  INV_X1    g318(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g319(.A(KEYINPUT37), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g320(.A1(new_n444_), .A2(new_n448_), .ZN(new_n458_));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n459_));
  NAND2_X1  g322(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g323(.A(new_n453_), .ZN(new_n461_));
  NAND3_X1  g324(.A1(new_n444_), .A2(new_n448_), .A3(KEYINPUT36), .ZN(new_n462_));
  NAND3_X1  g325(.A1(new_n460_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g326(.A(KEYINPUT37), .ZN(new_n464_));
  NAND3_X1  g327(.A1(new_n463_), .A2(new_n464_), .A3(new_n455_), .ZN(new_n465_));
  NAND2_X1  g328(.A1(new_n457_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g329(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g331(.A(new_n421_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g332(.A(new_n469_), .B(new_n388_), .ZN(new_n470_));
  XOR2_X1   g333(.A(G127gat), .B(G155gat), .Z(new_n471_));
  XNOR2_X1  g334(.A(new_n471_), .B(G211gat), .ZN(new_n472_));
  XOR2_X1   g335(.A(KEYINPUT16), .B(G183gat), .Z(new_n473_));
  XNOR2_X1  g336(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g337(.A1(new_n474_), .A2(KEYINPUT17), .ZN(new_n475_));
  NOR2_X1   g338(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g339(.A(new_n474_), .B(KEYINPUT17), .ZN(new_n477_));
  INV_X1    g340(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g341(.A(new_n476_), .B1(new_n470_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g342(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g343(.A1(new_n467_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g344(.A1(new_n438_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g345(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g346(.A1(new_n483_), .A2(new_n416_), .A3(new_n322_), .ZN(new_n484_));
  XNOR2_X1  g347(.A(new_n484_), .B(KEYINPUT38), .ZN(new_n485_));
  NAND2_X1  g348(.A1(new_n463_), .A2(new_n455_), .ZN(new_n486_));
  INV_X1    g349(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g350(.A1(new_n487_), .A2(new_n480_), .ZN(new_n488_));
  NAND2_X1  g351(.A1(new_n438_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g352(.A(new_n322_), .ZN(new_n490_));
  OAI21_X1  g353(.A(G1gat), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g354(.A1(new_n485_), .A2(new_n491_), .ZN(G1324gat));
  NOR2_X1   g355(.A1(new_n334_), .A2(new_n333_), .ZN(new_n493_));
  NAND3_X1  g356(.A1(new_n483_), .A2(new_n417_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g357(.A(KEYINPUT39), .ZN(new_n495_));
  NOR3_X1   g358(.A1(new_n437_), .A2(new_n487_), .A3(new_n480_), .ZN(new_n496_));
  NAND2_X1  g359(.A1(new_n496_), .A2(new_n493_), .ZN(new_n497_));
  AOI21_X1  g360(.A(new_n495_), .B1(new_n497_), .B2(G8gat), .ZN(new_n498_));
  AOI211_X1 g361(.A(KEYINPUT39), .B(new_n417_), .C1(new_n496_), .C2(new_n493_), .ZN(new_n499_));
  OAI21_X1  g362(.A(new_n494_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n501_));
  XNOR2_X1  g364(.A(new_n500_), .B(new_n501_), .ZN(G1325gat));
  INV_X1    g365(.A(G15gat), .ZN(new_n503_));
  AOI21_X1  g366(.A(new_n503_), .B1(new_n496_), .B2(new_n209_), .ZN(new_n504_));
  XNOR2_X1  g367(.A(new_n504_), .B(KEYINPUT41), .ZN(new_n505_));
  NAND3_X1  g368(.A1(new_n483_), .A2(new_n503_), .A3(new_n209_), .ZN(new_n506_));
  NAND2_X1  g369(.A1(new_n505_), .A2(new_n506_), .ZN(G1326gat));
  OAI21_X1  g370(.A(G22gat), .B1(new_n489_), .B2(new_n267_), .ZN(new_n508_));
  XNOR2_X1  g371(.A(new_n508_), .B(KEYINPUT42), .ZN(new_n509_));
  OR2_X1    g372(.A1(new_n267_), .A2(G22gat), .ZN(new_n510_));
  OAI21_X1  g373(.A(new_n509_), .B1(new_n482_), .B2(new_n510_), .ZN(G1327gat));
  INV_X1    g374(.A(KEYINPUT43), .ZN(new_n512_));
  AOI21_X1  g375(.A(new_n512_), .B1(new_n336_), .B2(new_n467_), .ZN(new_n513_));
  AOI211_X1 g376(.A(KEYINPUT43), .B(new_n466_), .C1(new_n330_), .C2(new_n335_), .ZN(new_n514_));
  OAI211_X1 g377(.A(new_n480_), .B(new_n436_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  INV_X1    g378(.A(KEYINPUT44), .ZN(new_n516_));
  NAND2_X1  g379(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI211_X1 g380(.A(new_n268_), .B(new_n331_), .C1(new_n323_), .C2(new_n328_), .ZN(new_n518_));
  NAND2_X1  g381(.A1(new_n304_), .A2(new_n305_), .ZN(new_n519_));
  NAND3_X1  g382(.A1(new_n325_), .A2(new_n299_), .A3(new_n327_), .ZN(new_n520_));
  OAI21_X1  g383(.A(new_n319_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g384(.A1(new_n521_), .A2(new_n267_), .ZN(new_n522_));
  AOI21_X1  g385(.A(new_n267_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n523_));
  NAND2_X1  g386(.A1(new_n523_), .A2(new_n490_), .ZN(new_n524_));
  NAND2_X1  g387(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g388(.A(new_n518_), .B1(new_n525_), .B2(new_n210_), .ZN(new_n526_));
  OAI21_X1  g389(.A(KEYINPUT43), .B1(new_n526_), .B2(new_n466_), .ZN(new_n527_));
  NAND3_X1  g390(.A1(new_n336_), .A2(new_n512_), .A3(new_n467_), .ZN(new_n528_));
  NAND2_X1  g391(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g392(.A1(new_n529_), .A2(KEYINPUT44), .A3(new_n480_), .A4(new_n436_), .ZN(new_n530_));
  NAND3_X1  g393(.A1(new_n517_), .A2(new_n322_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g394(.A1(new_n531_), .A2(G29gat), .ZN(new_n532_));
  NOR3_X1   g395(.A1(new_n437_), .A2(new_n486_), .A3(new_n479_), .ZN(new_n533_));
  INV_X1    g396(.A(new_n533_), .ZN(new_n534_));
  OR2_X1    g397(.A1(new_n490_), .A2(G29gat), .ZN(new_n535_));
  OAI21_X1  g398(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(G1328gat));
  NAND3_X1  g399(.A1(new_n517_), .A2(new_n493_), .A3(new_n530_), .ZN(new_n537_));
  NAND2_X1  g400(.A1(new_n537_), .A2(G36gat), .ZN(new_n538_));
  INV_X1    g401(.A(new_n493_), .ZN(new_n539_));
  NOR2_X1   g402(.A1(new_n539_), .A2(G36gat), .ZN(new_n540_));
  NAND2_X1  g403(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g404(.A(new_n541_), .B(KEYINPUT45), .ZN(new_n542_));
  NAND2_X1  g405(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g406(.A(KEYINPUT46), .ZN(new_n544_));
  NAND2_X1  g407(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g408(.A1(new_n538_), .A2(KEYINPUT46), .A3(new_n542_), .ZN(new_n546_));
  NAND2_X1  g409(.A1(new_n545_), .A2(new_n546_), .ZN(G1329gat));
  NAND3_X1  g410(.A1(new_n517_), .A2(new_n209_), .A3(new_n530_), .ZN(new_n548_));
  NAND2_X1  g411(.A1(new_n548_), .A2(G43gat), .ZN(new_n549_));
  OR3_X1    g412(.A1(new_n534_), .A2(G43gat), .A3(new_n210_), .ZN(new_n550_));
  NAND2_X1  g413(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g414(.A(KEYINPUT47), .ZN(new_n552_));
  NAND2_X1  g415(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g416(.A1(new_n549_), .A2(KEYINPUT47), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g417(.A1(new_n553_), .A2(new_n554_), .ZN(G1330gat));
  NAND3_X1  g418(.A1(new_n517_), .A2(new_n268_), .A3(new_n530_), .ZN(new_n556_));
  NAND2_X1  g419(.A1(new_n556_), .A2(G50gat), .ZN(new_n557_));
  OR2_X1    g420(.A1(new_n267_), .A2(G50gat), .ZN(new_n558_));
  OAI21_X1  g421(.A(new_n557_), .B1(new_n534_), .B2(new_n558_), .ZN(G1331gat));
  INV_X1    g422(.A(new_n435_), .ZN(new_n560_));
  INV_X1    g423(.A(new_n403_), .ZN(new_n561_));
  NOR3_X1   g424(.A1(new_n526_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AND2_X1   g425(.A1(new_n562_), .A2(new_n481_), .ZN(new_n563_));
  AOI21_X1  g426(.A(G57gat), .B1(new_n563_), .B2(new_n322_), .ZN(new_n564_));
  AND2_X1   g427(.A1(new_n562_), .A2(new_n488_), .ZN(new_n565_));
  AND2_X1   g428(.A1(new_n322_), .A2(G57gat), .ZN(new_n566_));
  AOI21_X1  g429(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(G1332gat));
  INV_X1    g430(.A(G64gat), .ZN(new_n568_));
  NAND3_X1  g431(.A1(new_n563_), .A2(new_n568_), .A3(new_n493_), .ZN(new_n569_));
  NAND2_X1  g432(.A1(new_n565_), .A2(new_n493_), .ZN(new_n570_));
  NAND2_X1  g433(.A1(new_n570_), .A2(G64gat), .ZN(new_n571_));
  AND2_X1   g434(.A1(new_n571_), .A2(KEYINPUT48), .ZN(new_n572_));
  NOR2_X1   g435(.A1(new_n571_), .A2(KEYINPUT48), .ZN(new_n573_));
  OAI21_X1  g436(.A(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(G1333gat));
  NAND3_X1  g437(.A1(new_n563_), .A2(new_n182_), .A3(new_n209_), .ZN(new_n575_));
  NAND2_X1  g438(.A1(new_n565_), .A2(new_n209_), .ZN(new_n576_));
  NAND2_X1  g439(.A1(new_n576_), .A2(G71gat), .ZN(new_n577_));
  AND2_X1   g440(.A1(new_n577_), .A2(KEYINPUT49), .ZN(new_n578_));
  NOR2_X1   g441(.A1(new_n577_), .A2(KEYINPUT49), .ZN(new_n579_));
  OAI21_X1  g442(.A(new_n575_), .B1(new_n578_), .B2(new_n579_), .ZN(G1334gat));
  INV_X1    g443(.A(G78gat), .ZN(new_n581_));
  NAND3_X1  g444(.A1(new_n563_), .A2(new_n581_), .A3(new_n268_), .ZN(new_n582_));
  NAND2_X1  g445(.A1(new_n565_), .A2(new_n268_), .ZN(new_n583_));
  NAND2_X1  g446(.A1(new_n583_), .A2(G78gat), .ZN(new_n584_));
  AND2_X1   g447(.A1(new_n584_), .A2(KEYINPUT50), .ZN(new_n585_));
  NOR2_X1   g448(.A1(new_n584_), .A2(KEYINPUT50), .ZN(new_n586_));
  OAI21_X1  g449(.A(new_n582_), .B1(new_n585_), .B2(new_n586_), .ZN(G1335gat));
  NOR2_X1   g450(.A1(new_n560_), .A2(new_n479_), .ZN(new_n588_));
  INV_X1    g451(.A(new_n588_), .ZN(new_n589_));
  NOR4_X1   g452(.A1(new_n526_), .A2(new_n486_), .A3(new_n561_), .A4(new_n589_), .ZN(new_n590_));
  AOI21_X1  g453(.A(G85gat), .B1(new_n590_), .B2(new_n322_), .ZN(new_n591_));
  AOI211_X1 g454(.A(new_n561_), .B(new_n589_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n592_));
  NOR2_X1   g455(.A1(new_n490_), .A2(new_n340_), .ZN(new_n593_));
  AOI21_X1  g456(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(G1336gat));
  AOI21_X1  g457(.A(G92gat), .B1(new_n590_), .B2(new_n493_), .ZN(new_n595_));
  NOR2_X1   g458(.A1(new_n539_), .A2(new_n341_), .ZN(new_n596_));
  AOI21_X1  g459(.A(new_n595_), .B1(new_n592_), .B2(new_n596_), .ZN(G1337gat));
  NAND4_X1  g460(.A1(new_n590_), .A2(new_n350_), .A3(new_n352_), .A4(new_n209_), .ZN(new_n598_));
  AND2_X1   g461(.A1(new_n592_), .A2(new_n209_), .ZN(new_n599_));
  OAI21_X1  g462(.A(new_n598_), .B1(new_n599_), .B2(new_n183_), .ZN(new_n600_));
  XNOR2_X1  g463(.A(new_n600_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g464(.A1(new_n590_), .A2(new_n351_), .A3(new_n268_), .ZN(new_n602_));
  NAND4_X1  g465(.A1(new_n529_), .A2(new_n268_), .A3(new_n403_), .A4(new_n588_), .ZN(new_n603_));
  INV_X1    g466(.A(KEYINPUT52), .ZN(new_n604_));
  AND3_X1   g467(.A1(new_n603_), .A2(new_n604_), .A3(G106gat), .ZN(new_n605_));
  AOI21_X1  g468(.A(new_n604_), .B1(new_n603_), .B2(G106gat), .ZN(new_n606_));
  OAI21_X1  g469(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g470(.A1(new_n607_), .A2(KEYINPUT53), .ZN(new_n608_));
  INV_X1    g471(.A(KEYINPUT53), .ZN(new_n609_));
  OAI211_X1 g472(.A(new_n609_), .B(new_n602_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g473(.A1(new_n608_), .A2(new_n610_), .ZN(G1339gat));
  NOR3_X1   g474(.A1(new_n493_), .A2(new_n490_), .A3(new_n210_), .ZN(new_n612_));
  INV_X1    g475(.A(new_n398_), .ZN(new_n613_));
  NOR2_X1   g476(.A1(new_n435_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g477(.A(KEYINPUT55), .ZN(new_n615_));
  NAND2_X1  g478(.A1(new_n390_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g479(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT55), .A4(new_n389_), .ZN(new_n617_));
  AND3_X1   g480(.A1(new_n379_), .A2(new_n389_), .A3(new_n374_), .ZN(new_n618_));
  OAI211_X1 g481(.A(new_n616_), .B(new_n617_), .C1(new_n337_), .C2(new_n618_), .ZN(new_n619_));
  AND3_X1   g482(.A1(new_n619_), .A2(KEYINPUT56), .A3(new_n396_), .ZN(new_n620_));
  AOI21_X1  g483(.A(KEYINPUT56), .B1(new_n619_), .B2(new_n396_), .ZN(new_n621_));
  OAI21_X1  g484(.A(new_n614_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g485(.A1(new_n426_), .A2(new_n423_), .ZN(new_n623_));
  NAND2_X1  g486(.A1(new_n422_), .A2(new_n424_), .ZN(new_n624_));
  OAI211_X1 g487(.A(new_n432_), .B(new_n623_), .C1(new_n624_), .C2(new_n423_), .ZN(new_n625_));
  AND2_X1   g488(.A1(new_n625_), .A2(new_n434_), .ZN(new_n626_));
  NAND2_X1  g489(.A1(new_n399_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g490(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g491(.A(KEYINPUT57), .B1(new_n628_), .B2(new_n486_), .ZN(new_n629_));
  INV_X1    g492(.A(KEYINPUT57), .ZN(new_n630_));
  AOI211_X1 g493(.A(new_n630_), .B(new_n487_), .C1(new_n622_), .C2(new_n627_), .ZN(new_n631_));
  NOR2_X1   g494(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g495(.A1(new_n626_), .A2(new_n398_), .ZN(new_n633_));
  OAI21_X1  g496(.A(new_n633_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n634_));
  INV_X1    g497(.A(KEYINPUT58), .ZN(new_n635_));
  NAND2_X1  g498(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g499(.A(KEYINPUT58), .B(new_n633_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n637_));
  NAND3_X1  g500(.A1(new_n636_), .A2(new_n467_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g501(.A(new_n479_), .B1(new_n632_), .B2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g502(.A1(new_n561_), .A2(new_n466_), .A3(new_n479_), .A4(new_n435_), .ZN(new_n640_));
  INV_X1    g503(.A(KEYINPUT54), .ZN(new_n641_));
  XNOR2_X1  g504(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  OAI211_X1 g505(.A(new_n267_), .B(new_n612_), .C1(new_n639_), .C2(new_n642_), .ZN(new_n643_));
  INV_X1    g506(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g507(.A(G113gat), .B1(new_n644_), .B2(new_n560_), .ZN(new_n645_));
  INV_X1    g508(.A(KEYINPUT59), .ZN(new_n646_));
  NAND2_X1  g509(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g510(.A1(new_n628_), .A2(new_n486_), .ZN(new_n648_));
  NAND2_X1  g511(.A1(new_n648_), .A2(new_n630_), .ZN(new_n649_));
  NAND3_X1  g512(.A1(new_n628_), .A2(KEYINPUT57), .A3(new_n486_), .ZN(new_n650_));
  NAND3_X1  g513(.A1(new_n649_), .A2(new_n650_), .A3(new_n638_), .ZN(new_n651_));
  NAND2_X1  g514(.A1(new_n651_), .A2(new_n480_), .ZN(new_n652_));
  INV_X1    g515(.A(new_n642_), .ZN(new_n653_));
  NAND2_X1  g516(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g517(.A1(new_n654_), .A2(KEYINPUT59), .A3(new_n267_), .A4(new_n612_), .ZN(new_n655_));
  AOI21_X1  g518(.A(new_n435_), .B1(new_n647_), .B2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g519(.A(new_n645_), .B1(new_n656_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g520(.A(new_n172_), .B1(new_n561_), .B2(KEYINPUT60), .ZN(new_n658_));
  OAI211_X1 g521(.A(new_n644_), .B(new_n658_), .C1(KEYINPUT60), .C2(new_n172_), .ZN(new_n659_));
  AOI21_X1  g522(.A(new_n561_), .B1(new_n647_), .B2(new_n655_), .ZN(new_n660_));
  OAI21_X1  g523(.A(new_n659_), .B1(new_n660_), .B2(new_n172_), .ZN(G1341gat));
  AOI21_X1  g524(.A(G127gat), .B1(new_n644_), .B2(new_n479_), .ZN(new_n662_));
  AOI21_X1  g525(.A(new_n480_), .B1(new_n647_), .B2(new_n655_), .ZN(new_n663_));
  AOI21_X1  g526(.A(new_n662_), .B1(new_n663_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g527(.A(G134gat), .B1(new_n644_), .B2(new_n487_), .ZN(new_n665_));
  AOI21_X1  g528(.A(new_n167_), .B1(new_n647_), .B2(new_n655_), .ZN(new_n666_));
  AOI21_X1  g529(.A(new_n665_), .B1(new_n666_), .B2(new_n467_), .ZN(G1343gat));
  NOR2_X1   g530(.A1(new_n490_), .A2(new_n209_), .ZN(new_n668_));
  NAND4_X1  g531(.A1(new_n654_), .A2(new_n523_), .A3(new_n560_), .A4(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g532(.A(new_n669_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g533(.A1(new_n654_), .A2(new_n523_), .A3(new_n403_), .A4(new_n668_), .ZN(new_n671_));
  XNOR2_X1  g534(.A(new_n671_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g535(.A1(new_n654_), .A2(new_n479_), .A3(new_n523_), .A4(new_n668_), .ZN(new_n673_));
  XNOR2_X1  g536(.A(KEYINPUT61), .B(G155gat), .ZN(new_n674_));
  XNOR2_X1  g537(.A(new_n673_), .B(new_n674_), .ZN(G1346gat));
  AND3_X1   g538(.A1(new_n654_), .A2(new_n523_), .A3(new_n668_), .ZN(new_n676_));
  NAND2_X1  g539(.A1(new_n676_), .A2(new_n487_), .ZN(new_n677_));
  INV_X1    g540(.A(G162gat), .ZN(new_n678_));
  NOR2_X1   g541(.A1(new_n466_), .A2(new_n678_), .ZN(new_n679_));
  AOI22_X1  g542(.A1(new_n677_), .A2(new_n678_), .B1(new_n676_), .B2(new_n679_), .ZN(G1347gat));
  AOI21_X1  g543(.A(new_n642_), .B1(new_n480_), .B2(new_n651_), .ZN(new_n681_));
  NOR2_X1   g544(.A1(new_n681_), .A2(new_n268_), .ZN(new_n682_));
  NOR2_X1   g545(.A1(new_n539_), .A2(new_n331_), .ZN(new_n683_));
  NAND3_X1  g546(.A1(new_n682_), .A2(new_n560_), .A3(new_n683_), .ZN(new_n684_));
  NAND3_X1  g547(.A1(new_n684_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n685_));
  INV_X1    g548(.A(KEYINPUT62), .ZN(new_n686_));
  INV_X1    g549(.A(new_n683_), .ZN(new_n687_));
  NOR4_X1   g550(.A1(new_n681_), .A2(new_n268_), .A3(new_n435_), .A4(new_n687_), .ZN(new_n688_));
  INV_X1    g551(.A(G169gat), .ZN(new_n689_));
  OAI21_X1  g552(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g553(.A1(new_n688_), .A2(new_n147_), .ZN(new_n691_));
  NAND3_X1  g554(.A1(new_n685_), .A2(new_n690_), .A3(new_n691_), .ZN(G1348gat));
  NAND3_X1  g555(.A1(new_n682_), .A2(new_n403_), .A3(new_n683_), .ZN(new_n693_));
  XNOR2_X1  g556(.A(new_n693_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g557(.A1(new_n654_), .A2(new_n479_), .A3(new_n267_), .A4(new_n683_), .ZN(new_n695_));
  AND2_X1   g558(.A1(new_n156_), .A2(new_n158_), .ZN(new_n696_));
  NOR2_X1   g559(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g560(.A(new_n697_), .B1(new_n138_), .B2(new_n695_), .ZN(G1350gat));
  NAND2_X1  g561(.A1(new_n682_), .A2(new_n683_), .ZN(new_n699_));
  OAI21_X1  g562(.A(G190gat), .B1(new_n699_), .B2(new_n466_), .ZN(new_n700_));
  NAND3_X1  g563(.A1(new_n487_), .A2(new_n159_), .A3(new_n161_), .ZN(new_n701_));
  OAI21_X1  g564(.A(new_n700_), .B1(new_n699_), .B2(new_n701_), .ZN(G1351gat));
  NOR3_X1   g565(.A1(new_n322_), .A2(new_n209_), .A3(new_n267_), .ZN(new_n703_));
  NAND4_X1  g566(.A1(new_n654_), .A2(new_n493_), .A3(new_n560_), .A4(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g567(.A(new_n704_), .B(G197gat), .ZN(G1352gat));
  AND3_X1   g568(.A1(new_n654_), .A2(new_n493_), .A3(new_n703_), .ZN(new_n706_));
  NAND2_X1  g569(.A1(new_n706_), .A2(new_n403_), .ZN(new_n707_));
  NAND2_X1  g570(.A1(new_n707_), .A2(G204gat), .ZN(new_n708_));
  NAND3_X1  g571(.A1(new_n706_), .A2(new_n216_), .A3(new_n403_), .ZN(new_n709_));
  NAND2_X1  g572(.A1(new_n708_), .A2(new_n709_), .ZN(G1353gat));
  NOR2_X1   g573(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n711_));
  AND2_X1   g574(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n712_));
  OAI211_X1 g575(.A(new_n706_), .B(new_n479_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n713_));
  AND2_X1   g576(.A1(new_n706_), .A2(new_n479_), .ZN(new_n714_));
  OAI21_X1  g577(.A(new_n713_), .B1(new_n714_), .B2(new_n711_), .ZN(G1354gat));
  NAND2_X1  g578(.A1(new_n706_), .A2(new_n487_), .ZN(new_n716_));
  INV_X1    g579(.A(G218gat), .ZN(new_n717_));
  NOR2_X1   g580(.A1(new_n466_), .A2(new_n717_), .ZN(new_n718_));
  AOI22_X1  g581(.A1(new_n716_), .A2(new_n717_), .B1(new_n706_), .B2(new_n718_), .ZN(G1355gat));
endmodule


