//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT90), .ZN(new_n203_));
  XOR2_X1   g002(.A(G127gat), .B(G134gat), .Z(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT91), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT91), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT31), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT89), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G227gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n212_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT86), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n216_), .B(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n220_), .B2(KEYINPUT23), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT83), .B(G190gat), .Z(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(G183gat), .B2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT88), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT22), .B(G169gat), .Z(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n223_), .A2(KEYINPUT88), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n224_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n225_), .A2(new_n226_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n222_), .A2(KEYINPUT26), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G190gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT84), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(KEYINPUT26), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243_));
  INV_X1    g042(.A(G183gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT82), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT25), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n242_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n235_), .B(new_n237_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n220_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT87), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n220_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n252_), .B(new_n254_), .C1(new_n250_), .C2(new_n217_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n233_), .B1(new_n249_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT30), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G71gat), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(G71gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n215_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n259_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n212_), .B(new_n213_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G15gat), .B(G43gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G99gat), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n261_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT94), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT3), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n272_), .A2(KEYINPUT2), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT95), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT95), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n277_), .A2(new_n283_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G155gat), .B(G162gat), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n278_), .B(KEYINPUT92), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n270_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295_));
  INV_X1    g094(.A(KEYINPUT97), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G197gat), .ZN(new_n298_));
  AOI211_X1 g097(.A(new_n294_), .B(new_n295_), .C1(new_n296_), .C2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G197gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G204gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n295_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT21), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(new_n302_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n293_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT96), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G78gat), .B(G106gat), .Z(new_n314_));
  NAND3_X1  g113(.A1(new_n293_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT98), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n318_));
  XOR2_X1   g117(.A(G22gat), .B(G50gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT28), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n318_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n313_), .A2(new_n315_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n314_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n316_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n322_), .A2(new_n326_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT18), .B(G64gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G92gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n257_), .B2(new_n308_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n244_), .A2(new_n240_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n230_), .B1(new_n255_), .B2(new_n338_), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n227_), .A2(KEYINPUT99), .A3(new_n234_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT99), .B1(new_n227_), .B2(new_n234_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n236_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AND4_X1   g144(.A1(new_n221_), .A2(new_n342_), .A3(new_n235_), .A4(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n307_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n347_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n308_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n233_), .B(new_n307_), .C1(new_n249_), .C2(new_n256_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n355_), .A2(KEYINPUT20), .A3(new_n351_), .A4(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n335_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(KEYINPUT101), .ZN(new_n360_));
  OR3_X1    g159(.A1(new_n339_), .A2(KEYINPUT101), .A3(new_n346_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n307_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n352_), .B1(new_n362_), .B2(new_n337_), .ZN(new_n363_));
  AND4_X1   g162(.A1(KEYINPUT20), .A2(new_n355_), .A3(new_n352_), .A4(new_n356_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n335_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(KEYINPUT27), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367_));
  INV_X1    g166(.A(new_n357_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n351_), .B1(new_n337_), .B2(new_n348_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n334_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n370_), .B2(new_n358_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n330_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n210_), .A2(new_n292_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n205_), .A2(new_n206_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n286_), .A2(new_n375_), .A3(new_n291_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT100), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT100), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n374_), .A2(new_n382_), .A3(KEYINPUT4), .A4(new_n376_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n210_), .A2(new_n292_), .A3(new_n378_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n379_), .A2(new_n381_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n377_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n380_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(G1gat), .B(G29gat), .Z(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n385_), .A2(new_n394_), .A3(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n269_), .A2(new_n373_), .A3(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT32), .B(new_n334_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n385_), .A2(new_n394_), .A3(new_n387_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n394_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n399_), .B(new_n401_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT102), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n370_), .A2(new_n358_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(KEYINPUT33), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n386_), .A2(new_n381_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n379_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n392_), .B(new_n409_), .C1(new_n410_), .C2(new_n381_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n395_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n407_), .A2(new_n408_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n396_), .A2(KEYINPUT102), .A3(new_n401_), .A4(new_n399_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n406_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n329_), .A2(new_n396_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n372_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n416_), .A2(new_n329_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n398_), .B1(new_n419_), .B2(new_n269_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT73), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT13), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n421_), .A2(KEYINPUT13), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G85gat), .A2(G92gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT9), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT64), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT10), .B(G99gat), .Z(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n425_), .A2(new_n427_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT9), .A3(new_n424_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(new_n439_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT10), .B(G99gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(G106gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT64), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n437_), .A3(KEYINPUT65), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT65), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT7), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT66), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n431_), .A2(new_n432_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n449_), .A2(new_n451_), .A3(new_n457_), .A4(new_n452_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT8), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n425_), .A2(new_n426_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n460_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n447_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n459_), .A2(new_n461_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT8), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT67), .A3(new_n447_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G57gat), .B(G64gat), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n474_));
  XOR2_X1   g273(.A(G71gat), .B(G78gat), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n474_), .A2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT68), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n466_), .A2(new_n471_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT69), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT69), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n447_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n478_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(KEYINPUT12), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G230gat), .A2(G233gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n479_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n464_), .A2(new_n465_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT67), .B1(new_n470_), .B2(new_n447_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n490_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n482_), .A2(new_n488_), .A3(new_n489_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT71), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT69), .B1(new_n462_), .B2(new_n463_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n468_), .A2(new_n484_), .A3(new_n469_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n478_), .B1(new_n499_), .B2(new_n447_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n466_), .A2(new_n471_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n500_), .A2(KEYINPUT12), .B1(new_n501_), .B2(new_n490_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n502_), .A2(KEYINPUT71), .A3(new_n489_), .A4(new_n482_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n493_), .A2(new_n480_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(G230gat), .A3(G233gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G120gat), .B(G148gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n297_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT5), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(new_n226_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n504_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(KEYINPUT72), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT72), .B1(new_n513_), .B2(new_n514_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n422_), .B(new_n423_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n517_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n519_), .A2(new_n515_), .A3(new_n421_), .A4(KEYINPUT13), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT81), .ZN(new_n522_));
  XOR2_X1   g321(.A(G15gat), .B(G22gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(G1gat), .A2(G8gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(KEYINPUT14), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT78), .ZN(new_n526_));
  XOR2_X1   g325(.A(G1gat), .B(G8gat), .Z(new_n527_));
  AND2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  INV_X1    g330(.A(G43gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G50gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n522_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n534_), .B(KEYINPUT15), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(new_n530_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(KEYINPUT81), .B2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n526_), .B(new_n527_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n534_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(new_n225_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n300_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n521_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT75), .B(G134gat), .ZN(new_n556_));
  INV_X1    g355(.A(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n486_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(new_n537_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n501_), .A2(new_n535_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT74), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(KEYINPUT35), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n569_), .A2(KEYINPUT35), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n564_), .A2(new_n571_), .A3(new_n572_), .A4(new_n565_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n562_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n562_), .A3(new_n573_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT77), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n576_), .A2(new_n581_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n578_), .A2(KEYINPUT76), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(KEYINPUT76), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n576_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT37), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n478_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n530_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n543_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT68), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT16), .B(G183gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(KEYINPUT79), .A3(KEYINPUT17), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT79), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n594_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT80), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AND4_X1   g408(.A1(new_n420_), .A2(new_n555_), .A3(new_n588_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n396_), .B(KEYINPUT103), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n611_), .A2(G1gat), .A3(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT38), .Z(new_n614_));
  AND2_X1   g413(.A1(new_n576_), .A2(new_n578_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n420_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT104), .B1(new_n420_), .B2(new_n616_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n607_), .B(new_n555_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n397_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(KEYINPUT105), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n625_));
  OAI211_X1 g424(.A(G8gat), .B(new_n625_), .C1(new_n621_), .C2(new_n418_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n617_), .B(new_n618_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n629_), .A2(new_n607_), .A3(new_n372_), .A4(new_n555_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n627_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(G8gat), .A3(new_n631_), .A4(new_n625_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n611_), .A2(G8gat), .A3(new_n418_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n628_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(new_n269_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G15gat), .B1(new_n621_), .B2(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT41), .ZN(new_n639_));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n610_), .A2(new_n640_), .A3(new_n269_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT107), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(KEYINPUT41), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT108), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n639_), .A2(new_n642_), .A3(new_n646_), .A4(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1326gat));
  OAI21_X1  g447(.A(G22gat), .B1(new_n621_), .B2(new_n329_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n329_), .A2(G22gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n611_), .B2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(new_n420_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n616_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n521_), .A2(new_n554_), .A3(new_n609_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n396_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n588_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(KEYINPUT109), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n420_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(KEYINPUT109), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n420_), .B2(new_n658_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n420_), .A2(new_n658_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n664_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n420_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n655_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n667_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n612_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n657_), .B1(new_n676_), .B2(G29gat), .ZN(G1328gat));
  AOI21_X1  g476(.A(KEYINPUT110), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n678_));
  OAI21_X1  g477(.A(G36gat), .B1(new_n675_), .B2(new_n418_), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n656_), .A2(new_n680_), .A3(new_n372_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT45), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n656_), .A2(new_n683_), .A3(new_n680_), .A4(new_n372_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n678_), .B1(new_n679_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(new_n685_), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT111), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1329gat));
  INV_X1    g490(.A(new_n656_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n532_), .B1(new_n692_), .B2(new_n637_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n269_), .A2(G43gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n675_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g495(.A(G50gat), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n675_), .A2(new_n697_), .A3(new_n329_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G50gat), .B1(new_n656_), .B2(new_n330_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1331gat));
  INV_X1    g499(.A(new_n521_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n554_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n703_), .A2(new_n420_), .A3(new_n588_), .A4(new_n609_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT112), .ZN(new_n705_));
  INV_X1    g504(.A(new_n612_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n629_), .A2(new_n609_), .A3(new_n703_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n397_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(G57gat), .B2(new_n709_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n708_), .B2(new_n418_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  INV_X1    g511(.A(new_n705_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n418_), .A2(G64gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n708_), .B2(new_n637_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n713_), .A2(G71gat), .A3(new_n637_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n708_), .B2(new_n329_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT114), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n720_), .B(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n329_), .A2(G78gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT115), .Z(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n713_), .B2(new_n725_), .ZN(G1335gat));
  NAND3_X1  g525(.A1(new_n521_), .A2(new_n554_), .A3(new_n608_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n727_), .A2(new_n728_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n666_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n396_), .A2(G85gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT117), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n653_), .A2(new_n727_), .A3(new_n616_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n706_), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n731_), .A2(new_n733_), .B1(new_n735_), .B2(G85gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT118), .ZN(G1336gat));
  AOI21_X1  g536(.A(G92gat), .B1(new_n734_), .B2(new_n372_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n731_), .A2(new_n418_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g539(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n734_), .A2(new_n436_), .A3(new_n269_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n666_), .A2(new_n269_), .A3(new_n729_), .A4(new_n730_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n743_), .A2(KEYINPUT119), .A3(G99gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT119), .B1(new_n743_), .B2(G99gat), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n741_), .B(new_n742_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n746_));
  OR2_X1    g545(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(G1338gat));
  NAND3_X1  g547(.A1(new_n734_), .A2(new_n437_), .A3(new_n330_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n666_), .A2(new_n330_), .A3(new_n729_), .A4(new_n730_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n608_), .A2(new_n702_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT121), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(new_n520_), .A3(new_n518_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n756_), .A2(KEYINPUT121), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n758_), .A2(new_n759_), .A3(new_n588_), .A4(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n757_), .A2(new_n588_), .A3(new_n520_), .A4(new_n518_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT54), .B1(new_n763_), .B2(new_n760_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT122), .B1(new_n504_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT122), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n770_), .B(KEYINPUT55), .C1(new_n496_), .C2(new_n503_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n494_), .A2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n502_), .A2(new_n482_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(G230gat), .A3(G233gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n769_), .A2(new_n771_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n767_), .B1(new_n776_), .B2(new_n511_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT123), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n504_), .A2(new_n768_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n770_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n775_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n504_), .A2(KEYINPUT122), .A3(new_n768_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n777_), .A2(new_n778_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n540_), .A2(new_n545_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n544_), .A2(new_n541_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n549_), .A3(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n551_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n514_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n766_), .B1(new_n785_), .B2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n512_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n790_), .B1(new_n794_), .B2(KEYINPUT123), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n777_), .A2(new_n778_), .A3(new_n784_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(KEYINPUT58), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n658_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT124), .ZN(new_n799_));
  INV_X1    g598(.A(new_n514_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n554_), .A2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n794_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n789_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n616_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n807_), .B(new_n615_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT124), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n793_), .A2(new_n810_), .A3(new_n658_), .A4(new_n797_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n799_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n607_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n765_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n706_), .A2(new_n269_), .A3(new_n373_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n702_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT59), .B1(new_n814_), .B2(new_n815_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n609_), .B1(new_n809_), .B2(new_n798_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n819_), .A2(new_n765_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n815_), .A2(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n702_), .A2(G113gat), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT125), .Z(new_n825_));
  AOI21_X1  g624(.A(new_n817_), .B1(new_n823_), .B2(new_n825_), .ZN(G1340gat));
  NAND3_X1  g625(.A1(new_n818_), .A2(new_n521_), .A3(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n701_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n816_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n814_), .A2(new_n815_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n608_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n818_), .A2(new_n822_), .A3(G127gat), .A4(new_n607_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1342gat));
  INV_X1    g636(.A(G134gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n834_), .B2(new_n616_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT126), .B(G134gat), .Z(new_n840_));
  NAND4_X1  g639(.A1(new_n818_), .A2(new_n822_), .A3(new_n658_), .A4(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n372_), .A2(new_n329_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n814_), .A2(new_n269_), .A3(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n702_), .A3(new_n706_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G141gat), .ZN(new_n847_));
  NOR4_X1   g646(.A1(new_n814_), .A2(new_n269_), .A3(new_n612_), .A4(new_n844_), .ZN(new_n848_));
  INV_X1    g647(.A(G141gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n702_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1344gat));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n521_), .A3(new_n706_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G148gat), .ZN(new_n853_));
  INV_X1    g652(.A(G148gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(new_n854_), .A3(new_n521_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1345gat));
  NAND2_X1  g655(.A1(new_n812_), .A2(new_n813_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n765_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n269_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n859_), .A2(new_n706_), .A3(new_n609_), .A4(new_n843_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n845_), .A2(new_n706_), .A3(new_n609_), .A4(new_n861_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1346gat));
  NAND2_X1  g664(.A1(new_n848_), .A2(new_n615_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n588_), .A2(new_n557_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT127), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n866_), .A2(new_n557_), .B1(new_n848_), .B2(new_n868_), .ZN(G1347gat));
  NOR3_X1   g668(.A1(new_n637_), .A2(new_n706_), .A3(new_n418_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n329_), .B(new_n870_), .C1(new_n819_), .C2(new_n765_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n871_), .A2(new_n554_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n871_), .B2(new_n554_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n873_), .B(new_n876_), .C1(new_n229_), .C2(new_n872_), .ZN(G1348gat));
  NOR4_X1   g676(.A1(new_n814_), .A2(new_n226_), .A3(new_n330_), .A4(new_n701_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n871_), .A2(new_n701_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n870_), .A2(new_n878_), .B1(new_n879_), .B2(new_n226_), .ZN(G1349gat));
  NOR3_X1   g679(.A1(new_n871_), .A2(new_n813_), .A3(new_n343_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n814_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n882_), .A2(new_n329_), .A3(new_n609_), .A4(new_n870_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n883_), .B2(new_n244_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n871_), .B2(new_n588_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n615_), .A2(new_n344_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n871_), .B2(new_n886_), .ZN(G1351gat));
  NAND2_X1  g686(.A1(new_n417_), .A2(new_n372_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n859_), .A2(new_n702_), .A3(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g690(.A1(new_n859_), .A2(new_n521_), .A3(new_n889_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g692(.A(KEYINPUT63), .B(G211gat), .Z(new_n894_));
  AND4_X1   g693(.A1(new_n607_), .A2(new_n859_), .A3(new_n889_), .A4(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n859_), .A2(new_n607_), .A3(new_n889_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n859_), .A2(new_n615_), .A3(new_n889_), .ZN(new_n900_));
  NOR4_X1   g699(.A1(new_n814_), .A2(new_n899_), .A3(new_n269_), .A4(new_n888_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n658_), .ZN(G1355gat));
endmodule


