//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT88), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n204_), .A2(KEYINPUT1), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G155gat), .ZN(new_n207_));
  INV_X1    g006(.A(G162gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT1), .B1(new_n204_), .B2(new_n205_), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n210_), .A2(KEYINPUT89), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(KEYINPUT89), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n209_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G141gat), .ZN(new_n219_));
  INV_X1    g018(.A(G148gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT3), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n214_), .A2(KEYINPUT90), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT2), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n214_), .A2(KEYINPUT90), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT91), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT91), .A4(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n204_), .A2(new_n205_), .B1(G155gat), .B2(G162gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT92), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT92), .ZN(new_n237_));
  AOI211_X1 g036(.A(new_n237_), .B(new_n234_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n218_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n239_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT28), .B1(new_n239_), .B2(KEYINPUT29), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G22gat), .B(G50gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246_));
  INV_X1    g045(.A(new_n217_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n210_), .B(KEYINPUT89), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n209_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(G141gat), .B2(G148gat), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n227_), .A2(new_n251_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT91), .B1(new_n252_), .B2(new_n226_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n232_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n235_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n237_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n233_), .A2(KEYINPUT92), .A3(new_n235_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n249_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n246_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n245_), .B1(new_n240_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n244_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G197gat), .B(G204gat), .Z(new_n263_));
  OR2_X1    g062(.A1(new_n263_), .A2(KEYINPUT21), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(KEYINPUT21), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n265_), .A2(new_n266_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT93), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G228gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n273_), .A3(new_n271_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G78gat), .B(G106gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n262_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n276_), .B2(new_n271_), .ZN(new_n285_));
  AOI211_X1 g084(.A(new_n274_), .B(new_n270_), .C1(new_n239_), .C2(KEYINPUT29), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT94), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT94), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n275_), .A2(new_n277_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n289_), .A3(new_n278_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT95), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT95), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n287_), .A2(new_n289_), .A3(new_n292_), .A4(new_n278_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n280_), .A2(new_n244_), .A3(new_n261_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AND4_X1   g094(.A1(new_n284_), .A2(new_n291_), .A3(new_n293_), .A4(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n290_), .B2(KEYINPUT95), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n284_), .B1(new_n297_), .B2(new_n293_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n283_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT97), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT97), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n301_), .B(new_n283_), .C1(new_n296_), .C2(new_n298_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NAND3_X1  g105(.A1(new_n239_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT100), .Z(new_n309_));
  INV_X1    g108(.A(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n258_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n239_), .A2(new_n306_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n307_), .B(new_n309_), .C1(new_n313_), .C2(new_n303_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n309_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G85gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G57gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  AND3_X1   g118(.A1(new_n314_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n269_), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT24), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT78), .B(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT26), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n329_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT79), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(KEYINPUT80), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(KEYINPUT23), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n328_), .A2(new_n327_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(KEYINPUT81), .A3(new_n341_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n336_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n339_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n347_), .A2(KEYINPUT84), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n331_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n347_), .A2(new_n348_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT84), .B1(new_n337_), .B2(KEYINPUT23), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n349_), .B(new_n351_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n355_));
  AOI21_X1  g154(.A(G176gat), .B1(new_n355_), .B2(KEYINPUT82), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT22), .B(G169gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(KEYINPUT82), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT83), .ZN(new_n359_));
  INV_X1    g158(.A(new_n326_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n323_), .B1(new_n346_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n340_), .B1(G183gat), .B2(G190gat), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n326_), .A2(KEYINPUT98), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n326_), .A2(KEYINPUT98), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n364_), .A2(new_n365_), .B1(new_n325_), .B2(new_n357_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n349_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n329_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n334_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n341_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n367_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT20), .B1(new_n373_), .B2(new_n269_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n362_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n346_), .A2(new_n361_), .A3(new_n323_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n373_), .B2(new_n269_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n377_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT18), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT32), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n377_), .B1(new_n362_), .B2(new_n374_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n380_), .A2(new_n382_), .A3(new_n378_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n395_), .A2(new_n391_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n322_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT101), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n320_), .A2(KEYINPUT33), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n379_), .A2(new_n390_), .A3(new_n384_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n362_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n378_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n389_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n404_), .A3(KEYINPUT99), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT99), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n385_), .A2(new_n406_), .A3(new_n389_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n320_), .A2(KEYINPUT33), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n311_), .A2(new_n312_), .A3(new_n309_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n319_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n307_), .B1(new_n313_), .B2(new_n303_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n410_), .B(new_n411_), .C1(new_n412_), .C2(new_n309_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n400_), .A2(new_n408_), .A3(new_n409_), .A4(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT101), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n322_), .A2(new_n415_), .A3(new_n397_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n399_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n300_), .A2(new_n302_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n300_), .A2(new_n417_), .A3(KEYINPUT102), .A4(new_n302_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n300_), .A2(new_n302_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n322_), .A2(KEYINPUT103), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n322_), .A2(KEYINPUT103), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n408_), .A2(KEYINPUT27), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n395_), .A2(new_n389_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n401_), .A3(KEYINPUT27), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n420_), .A2(new_n421_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n346_), .A2(new_n361_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n435_), .A2(KEYINPUT86), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  INV_X1    g236(.A(G43gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT85), .B(G15gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n435_), .B2(KEYINPUT86), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n436_), .B(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n306_), .A2(KEYINPUT31), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n306_), .A2(KEYINPUT31), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n446_), .A2(KEYINPUT87), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n445_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n432_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n429_), .A2(KEYINPUT104), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT104), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n426_), .A2(new_n452_), .A3(new_n428_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n449_), .A2(new_n425_), .ZN(new_n455_));
  AND4_X1   g254(.A1(new_n300_), .A2(new_n454_), .A3(new_n302_), .A4(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n450_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G15gat), .B(G22gat), .Z(new_n459_));
  NAND2_X1  g258(.A1(G1gat), .A2(G8gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(KEYINPUT14), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT75), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G1gat), .B(G8gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(KEYINPUT15), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n474_), .A2(KEYINPUT77), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(KEYINPUT77), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n464_), .B(new_n467_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n473_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n475_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G113gat), .B(G141gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G169gat), .B(G197gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n483_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n458_), .A2(KEYINPUT105), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT105), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n456_), .B1(new_n432_), .B2(new_n449_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n486_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT13), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G85gat), .B(G92gat), .ZN(new_n494_));
  INV_X1    g293(.A(G92gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(KEYINPUT9), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(KEYINPUT9), .B2(new_n494_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT64), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT6), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT6), .B1(new_n500_), .B2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT65), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n494_), .A2(KEYINPUT8), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n501_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT7), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(KEYINPUT66), .B2(new_n504_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n504_), .A2(KEYINPUT66), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n494_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n522_));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n509_), .A2(new_n526_), .A3(new_n518_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(KEYINPUT12), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n519_), .A2(new_n531_), .A3(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G230gat), .A2(G233gat), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n528_), .A2(new_n529_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G230gat), .A3(G233gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(G120gat), .B(G148gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n538_), .A2(new_n540_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n493_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n538_), .A2(new_n540_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n545_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT13), .A3(new_n546_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n526_), .B(new_n555_), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n464_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT17), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n562_), .B(KEYINPUT17), .Z(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT69), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT36), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT71), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n467_), .ZN(new_n579_));
  OAI22_X1  g378(.A1(new_n519_), .A2(new_n579_), .B1(KEYINPUT35), .B2(new_n575_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n470_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n580_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n573_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT72), .ZN(new_n586_));
  INV_X1    g385(.A(new_n584_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n571_), .A2(KEYINPUT36), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT70), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n582_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n585_), .A2(KEYINPUT72), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT37), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n585_), .A2(new_n590_), .A3(KEYINPUT74), .A4(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n567_), .B1(new_n593_), .B2(new_n599_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n492_), .A2(new_n554_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(G1gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n425_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n585_), .A2(new_n590_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n489_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(new_n486_), .A3(new_n554_), .A4(new_n566_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n425_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n603_), .A2(new_n604_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n605_), .A2(new_n610_), .A3(new_n611_), .ZN(G1324gat));
  OAI21_X1  g411(.A(G8gat), .B1(new_n608_), .B2(new_n454_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT39), .ZN(new_n614_));
  INV_X1    g413(.A(G8gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n454_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n601_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(KEYINPUT40), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n608_), .B2(new_n449_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT41), .Z(new_n624_));
  INV_X1    g423(.A(G15gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n449_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n601_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(G1326gat));
  INV_X1    g427(.A(new_n422_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G22gat), .B1(new_n608_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n601_), .A2(new_n632_), .A3(new_n422_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n631_), .A2(KEYINPUT106), .A3(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1327gat));
  NAND4_X1  g437(.A1(new_n549_), .A2(new_n553_), .A3(new_n486_), .A4(new_n567_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT107), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n593_), .A2(new_n599_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n458_), .B2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n489_), .A2(KEYINPUT43), .A3(new_n643_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT44), .B(new_n641_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT108), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n489_), .B2(new_n643_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n418_), .A2(new_n419_), .B1(new_n422_), .B2(new_n430_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n626_), .B1(new_n650_), .B2(new_n421_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n642_), .B(new_n644_), .C1(new_n651_), .C2(new_n456_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n640_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT108), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n641_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n425_), .A3(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT109), .A3(G29gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT109), .B1(new_n660_), .B2(G29gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n606_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n566_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n554_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n609_), .A2(G29gat), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT110), .Z(new_n669_));
  OAI22_X1  g468(.A1(new_n661_), .A2(new_n662_), .B1(new_n667_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT111), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(KEYINPUT111), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n454_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n656_), .B2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n454_), .A2(G36gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT45), .B1(new_n666_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n666_), .A2(KEYINPUT45), .A3(new_n677_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n672_), .B(new_n673_), .C1(new_n676_), .C2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n653_), .A2(new_n654_), .A3(KEYINPUT44), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n654_), .B1(new_n653_), .B2(KEYINPUT44), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n675_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n679_), .A2(new_n680_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(KEYINPUT111), .A4(new_n671_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n682_), .A2(new_n688_), .ZN(G1329gat));
  NAND4_X1  g488(.A1(new_n656_), .A2(G43gat), .A3(new_n626_), .A4(new_n659_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n438_), .B1(new_n667_), .B2(new_n449_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(KEYINPUT47), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT47), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1330gat));
  INV_X1    g493(.A(G50gat), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n648_), .A2(new_n655_), .B1(new_n658_), .B2(new_n657_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n422_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n422_), .A2(new_n695_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT112), .Z(new_n699_));
  NOR2_X1   g498(.A1(new_n667_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT113), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n656_), .A2(new_n422_), .A3(new_n659_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G50gat), .ZN(new_n703_));
  INV_X1    g502(.A(new_n700_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT113), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n701_), .A2(new_n706_), .ZN(G1331gat));
  NAND2_X1  g506(.A1(new_n549_), .A2(new_n553_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n607_), .A2(new_n490_), .A3(new_n708_), .A4(new_n566_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n609_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n458_), .A2(new_n490_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(KEYINPUT114), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n554_), .B1(new_n711_), .B2(KEYINPUT114), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n600_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n609_), .A2(G57gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n710_), .B1(new_n715_), .B2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n709_), .B2(new_n454_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n454_), .A2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n715_), .B2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n709_), .B2(new_n449_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n449_), .A2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n715_), .B2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n709_), .B2(new_n629_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n629_), .A2(G78gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n715_), .B2(new_n728_), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n486_), .A2(new_n566_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n708_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT115), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n609_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n712_), .A2(new_n664_), .A3(new_n713_), .ZN(new_n736_));
  INV_X1    g535(.A(G85gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n425_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT116), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n734_), .B2(new_n454_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n616_), .A2(new_n495_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n736_), .B2(new_n742_), .ZN(G1337gat));
  NAND2_X1  g542(.A1(new_n733_), .A2(new_n626_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n744_), .A2(KEYINPUT117), .A3(G99gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT117), .B1(new_n744_), .B2(G99gat), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n626_), .A2(new_n506_), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n745_), .A2(new_n746_), .B1(new_n736_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g548(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n629_), .B(new_n732_), .C1(new_n649_), .C2(new_n652_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT118), .B1(new_n752_), .B2(new_n501_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n754_), .B(G106gat), .C1(new_n734_), .C2(new_n629_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n755_), .A3(KEYINPUT52), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n714_), .A2(new_n501_), .A3(new_n422_), .A4(new_n664_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(new_n753_), .B2(new_n755_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n759_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(new_n757_), .A3(new_n756_), .A4(new_n750_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT122), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n606_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n546_), .A2(new_n486_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n533_), .A2(new_n535_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n533_), .A2(KEYINPUT55), .A3(new_n535_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n538_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n773_), .B2(new_n545_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n533_), .A2(new_n535_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT67), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n772_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n770_), .A3(new_n769_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n551_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n767_), .B1(new_n774_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n482_), .B1(new_n477_), .B2(new_n472_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n472_), .B2(new_n471_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n484_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n552_), .B2(new_n546_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n766_), .B1(new_n781_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n764_), .A2(new_n765_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n766_), .B(new_n788_), .C1(new_n781_), .C2(new_n786_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n784_), .A2(new_n546_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n551_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(KEYINPUT121), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n774_), .A2(new_n796_), .A3(new_n780_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT58), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n643_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n567_), .B1(new_n792_), .B2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n554_), .A2(KEYINPUT120), .A3(new_n490_), .A4(new_n600_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n600_), .A2(new_n490_), .A3(new_n549_), .A4(new_n553_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n807_), .A3(KEYINPUT54), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n609_), .B1(new_n803_), .B2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n616_), .A2(new_n422_), .A3(new_n449_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n486_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n813_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n490_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n816_), .B1(new_n821_), .B2(new_n815_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n554_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n814_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n554_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1341gat));
  NAND2_X1  g626(.A1(new_n814_), .A2(new_n566_), .ZN(new_n828_));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT123), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT123), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n817_), .A2(new_n820_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n567_), .A2(new_n829_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n831_), .A2(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n814_), .A2(new_n837_), .A3(new_n606_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n643_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1343gat));
  NAND2_X1  g639(.A1(new_n422_), .A2(new_n449_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n616_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n790_), .A2(new_n791_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n799_), .A2(new_n801_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n644_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n566_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n808_), .A2(new_n810_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n425_), .B(new_n842_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n812_), .A2(KEYINPUT124), .A3(new_n842_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n490_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n219_), .ZN(G1344gat));
  AOI21_X1  g652(.A(new_n554_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(new_n220_), .ZN(G1345gat));
  AOI21_X1  g654(.A(new_n567_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT61), .B(G155gat), .Z(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  AOI211_X1 g657(.A(new_n208_), .B(new_n643_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n663_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT125), .B1(new_n860_), .B2(G162gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n803_), .A2(new_n811_), .ZN(new_n862_));
  AND4_X1   g661(.A1(KEYINPUT124), .A2(new_n862_), .A3(new_n425_), .A4(new_n842_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT124), .B1(new_n812_), .B2(new_n842_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n606_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n208_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n859_), .B1(new_n861_), .B2(new_n867_), .ZN(G1347gat));
  NAND2_X1  g667(.A1(new_n616_), .A2(new_n609_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n869_), .A2(new_n449_), .A3(new_n422_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n324_), .B1(new_n872_), .B2(new_n486_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n873_), .A2(KEYINPUT62), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n357_), .A3(new_n486_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(KEYINPUT62), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .ZN(G1348gat));
  NOR2_X1   g676(.A1(new_n871_), .A2(new_n554_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n325_), .ZN(G1349gat));
  NOR2_X1   g678(.A1(new_n871_), .A2(new_n567_), .ZN(new_n880_));
  MUX2_X1   g679(.A(G183gat), .B(new_n334_), .S(new_n880_), .Z(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n871_), .B2(new_n643_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n606_), .A2(new_n370_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n871_), .B2(new_n883_), .ZN(G1351gat));
  NOR2_X1   g683(.A1(new_n869_), .A2(new_n841_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n862_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n486_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g688(.A1(new_n886_), .A2(new_n554_), .ZN(new_n890_));
  AND2_X1   g689(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n890_), .B2(new_n892_), .ZN(G1353gat));
  NAND2_X1  g693(.A1(new_n887_), .A2(new_n566_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  AND2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n895_), .B2(new_n896_), .ZN(G1354gat));
  INV_X1    g698(.A(G218gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n887_), .A2(new_n900_), .A3(new_n606_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n886_), .A2(new_n643_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT127), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n901_), .B(new_n905_), .C1(new_n900_), .C2(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1355gat));
endmodule


