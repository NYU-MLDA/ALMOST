//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  AOI21_X1  g003(.A(KEYINPUT87), .B1(new_n204_), .B2(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  AOI22_X1  g007(.A1(new_n206_), .A2(new_n207_), .B1(new_n208_), .B2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n204_), .A2(G197gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(G204gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(new_n211_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n218_));
  INV_X1    g017(.A(new_n207_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n215_), .B(new_n218_), .C1(new_n219_), .C2(new_n205_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT89), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT89), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n217_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n213_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n235_));
  NAND3_X1  g034(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G141gat), .A2(G148gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n229_), .B(new_n231_), .C1(new_n240_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n241_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n234_), .A2(new_n236_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(G155gat), .A3(G162gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT83), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n227_), .B(new_n228_), .C1(new_n230_), .C2(new_n247_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n245_), .B(new_n246_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n226_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n203_), .B1(new_n225_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n244_), .A2(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT29), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n224_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n223_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n260_), .A3(new_n202_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G78gat), .B(G106gat), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT91), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n266_));
  INV_X1    g065(.A(G22gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G50gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n244_), .A2(new_n252_), .A3(KEYINPUT85), .A4(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(new_n274_), .A3(new_n270_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n254_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n263_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n265_), .A2(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n277_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(new_n275_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n281_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT91), .A4(new_n279_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT31), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT77), .B(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT25), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT78), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n296_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT79), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G183gat), .ZN(new_n310_));
  INV_X1    g109(.A(G190gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT23), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n306_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n295_), .A2(new_n299_), .A3(new_n305_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n307_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n291_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(G190gat), .ZN(new_n318_));
  OR2_X1    g117(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n302_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n315_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n315_), .B2(new_n324_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n289_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G120gat), .ZN(new_n330_));
  INV_X1    g129(.A(G127gat), .ZN(new_n331_));
  INV_X1    g130(.A(G134gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G113gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G127gat), .A2(G134gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n330_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(G120gat), .A3(new_n336_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G71gat), .B(G99gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT30), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n328_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n289_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n326_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n329_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n329_), .B2(new_n354_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n287_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(G1gat), .B(G29gat), .Z(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n255_), .A2(new_n342_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT98), .B1(new_n365_), .B2(KEYINPUT4), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n244_), .A2(new_n252_), .A3(new_n341_), .A4(new_n339_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(KEYINPUT4), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT98), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n255_), .A2(new_n369_), .A3(new_n370_), .A4(new_n342_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n376_));
  OAI211_X1 g175(.A(KEYINPUT33), .B(new_n364_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT33), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n363_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT18), .B(G64gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G92gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G8gat), .B(G36gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n303_), .A2(KEYINPUT94), .A3(new_n298_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT94), .B1(new_n303_), .B2(new_n298_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n301_), .A3(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(KEYINPUT25), .B(G183gat), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n290_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n296_), .A2(new_n298_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n316_), .A2(KEYINPUT95), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT95), .B1(new_n316_), .B2(new_n393_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n389_), .B(new_n392_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n314_), .B1(G183gat), .B2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n321_), .A2(KEYINPUT96), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n319_), .A2(new_n401_), .A3(new_n320_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n303_), .B1(new_n403_), .B2(new_n322_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n314_), .B(KEYINPUT97), .C1(G183gat), .C2(G190gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n225_), .A2(new_n396_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT92), .Z(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT19), .Z(new_n410_));
  NAND2_X1  g209(.A1(new_n315_), .A2(new_n324_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n260_), .A2(new_n411_), .ZN(new_n412_));
  AND4_X1   g211(.A1(KEYINPUT20), .A2(new_n407_), .A3(new_n410_), .A4(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n410_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n411_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT93), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n406_), .A2(new_n396_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n260_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n260_), .C2(new_n411_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI211_X1 g220(.A(new_n386_), .B(new_n413_), .C1(new_n414_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n414_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n413_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n385_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n366_), .A2(new_n368_), .A3(new_n373_), .A4(new_n371_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n365_), .A2(new_n374_), .A3(new_n367_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n363_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n381_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n379_), .B(new_n363_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n413_), .B1(new_n421_), .B2(new_n414_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT99), .A3(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n417_), .A2(new_n410_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n407_), .A2(KEYINPUT20), .A3(new_n412_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n414_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT99), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n431_), .B(new_n434_), .C1(new_n440_), .C2(new_n433_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n359_), .B1(new_n430_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n379_), .B(new_n364_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n282_), .A2(new_n286_), .A3(new_n357_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n357_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT27), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n432_), .A2(new_n385_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n438_), .A2(new_n386_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(KEYINPUT27), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n442_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G71gat), .B(G78gat), .Z(new_n455_));
  OR2_X1    g254(.A1(G57gat), .A2(G64gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n458_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(KEYINPUT11), .ZN(new_n463_));
  AND2_X1   g262(.A1(G57gat), .A2(G64gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G57gat), .A2(G64gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n461_), .B(KEYINPUT11), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n460_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT11), .B1(new_n464_), .B2(new_n465_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT66), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(new_n459_), .A3(new_n455_), .A4(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G1gat), .A2(G8gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT14), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G15gat), .A2(G22gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(G15gat), .A2(G22gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n473_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n483_), .A2(new_n473_), .A3(new_n480_), .A4(new_n474_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n472_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G231gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT72), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT16), .B(G183gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G211gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G127gat), .B(G155gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT17), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n489_), .B(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n488_), .A2(KEYINPUT17), .A3(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT34), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT35), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT69), .Z(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n516_), .A2(KEYINPUT65), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT8), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT10), .B(G99gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT64), .B(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n511_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n516_), .A2(KEYINPUT9), .A3(new_n517_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n517_), .A2(KEYINPUT9), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n520_), .A2(new_n522_), .B1(new_n525_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n269_), .A2(G43gat), .ZN(new_n533_));
  INV_X1    g332(.A(G43gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(G50gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G36gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G29gat), .ZN(new_n538_));
  INV_X1    g337(.A(G29gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G36gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n533_), .A2(new_n535_), .A3(new_n538_), .A4(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n532_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT70), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n533_), .A2(new_n535_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT15), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI22_X1  g352(.A1(new_n532_), .A2(new_n553_), .B1(KEYINPUT35), .B2(new_n502_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT70), .B1(new_n532_), .B2(new_n544_), .ZN(new_n555_));
  OR4_X1    g354(.A1(new_n504_), .A2(new_n547_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G190gat), .B(G218gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G134gat), .ZN(new_n558_));
  INV_X1    g357(.A(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n545_), .B(new_n546_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n504_), .B1(new_n561_), .B2(new_n554_), .ZN(new_n562_));
  AND4_X1   g361(.A1(new_n500_), .A2(new_n556_), .A3(new_n560_), .A4(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n560_), .B(new_n500_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n499_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NOR4_X1   g367(.A1(new_n563_), .A2(new_n565_), .A3(new_n567_), .A4(new_n499_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n454_), .A2(new_n498_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n532_), .A2(new_n472_), .B1(KEYINPUT67), .B2(KEYINPUT12), .ZN(new_n574_));
  NOR2_X1   g373(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n532_), .A2(new_n472_), .A3(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n468_), .A2(new_n471_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n525_), .A2(new_n528_), .A3(new_n530_), .A4(new_n529_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n513_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n521_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n575_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n573_), .B(new_n574_), .C1(new_n577_), .C2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n582_), .B(new_n472_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n573_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G120gat), .B(G148gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n586_), .B(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT13), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT73), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT73), .B1(new_n542_), .B2(new_n543_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n485_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n482_), .A2(new_n484_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n551_), .A2(new_n600_), .A3(new_n552_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(new_n599_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n485_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n544_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n542_), .A2(new_n543_), .A3(KEYINPUT73), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n600_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n604_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT75), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n334_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT75), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n612_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(G113gat), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(G113gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n334_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(G141gat), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT74), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n598_), .A2(new_n601_), .A3(new_n623_), .A4(new_n599_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n603_), .A2(new_n610_), .A3(new_n622_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n626_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n603_), .A2(new_n610_), .A3(new_n624_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n622_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n627_), .A2(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n595_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n572_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n478_), .A3(new_n431_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT38), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n563_), .A2(new_n565_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT100), .B1(new_n454_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n639_), .B(new_n566_), .C1(new_n442_), .C2(new_n453_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n497_), .A3(new_n632_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n443_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n636_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n636_), .A2(KEYINPUT101), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1324gat));
  NAND4_X1  g447(.A1(new_n641_), .A2(new_n497_), .A3(new_n452_), .A4(new_n632_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n649_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n633_), .A2(G8gat), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT102), .A3(new_n452_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT102), .B1(new_n654_), .B2(new_n452_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n652_), .B(new_n653_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  INV_X1    g458(.A(new_n357_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n633_), .A2(G15gat), .A3(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n642_), .A2(new_n660_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT41), .B1(new_n662_), .B2(G15gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(new_n287_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G22gat), .B1(new_n642_), .B2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT103), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT103), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n634_), .A2(new_n267_), .A3(new_n287_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n670_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .ZN(G1327gat));
  NOR2_X1   g473(.A1(new_n454_), .A2(new_n566_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n595_), .A2(new_n497_), .A3(new_n631_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n431_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT37), .B1(new_n637_), .B2(KEYINPUT71), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n569_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n430_), .A2(new_n441_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n358_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n448_), .A2(new_n451_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n287_), .A2(new_n660_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n282_), .A2(new_n357_), .A3(new_n286_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n431_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n681_), .B1(new_n683_), .B2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n571_), .B1(new_n442_), .B2(new_n453_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n690_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(KEYINPUT105), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n695_), .A2(new_n676_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n689_), .B2(KEYINPUT104), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n692_), .A2(new_n693_), .A3(new_n691_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n701_), .A2(new_n676_), .A3(new_n699_), .A4(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n697_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n443_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n679_), .B1(new_n705_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n678_), .A2(new_n537_), .A3(new_n452_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n684_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n537_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n708_), .B(KEYINPUT46), .C1(new_n709_), .C2(new_n537_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  AND2_X1   g513(.A1(new_n703_), .A2(new_n697_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n703_), .A2(new_n697_), .ZN(new_n716_));
  OAI211_X1 g515(.A(G43gat), .B(new_n357_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G43gat), .B1(new_n678_), .B2(new_n357_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n287_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G50gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n678_), .A2(new_n269_), .A3(new_n287_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n666_), .B1(new_n700_), .B2(new_n704_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n722_), .B(new_n725_), .C1(new_n727_), .C2(new_n269_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n595_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n625_), .B(new_n626_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n629_), .A2(new_n630_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n572_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n431_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n731_), .A2(new_n498_), .A3(new_n734_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n423_), .A2(new_n439_), .A3(new_n424_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n438_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n433_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n443_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n429_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n422_), .A2(new_n425_), .A3(new_n744_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n743_), .A2(new_n434_), .B1(new_n745_), .B2(new_n381_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n688_), .B1(new_n746_), .B2(new_n359_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n639_), .B1(new_n747_), .B2(new_n566_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n640_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n739_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n641_), .A2(KEYINPUT107), .A3(new_n739_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n431_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n738_), .B1(new_n754_), .B2(G57gat), .ZN(G1332gat));
  NOR2_X1   g554(.A1(new_n684_), .A2(G64gat), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT109), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n737_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n752_), .A2(new_n452_), .A3(new_n753_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G64gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT108), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(G64gat), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n761_), .A2(KEYINPUT48), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT48), .B1(new_n761_), .B2(new_n763_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n758_), .B1(new_n764_), .B2(new_n765_), .ZN(G1333gat));
  OR3_X1    g565(.A1(new_n736_), .A2(G71gat), .A3(new_n660_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n752_), .A2(new_n357_), .A3(new_n753_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G71gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1334gat));
  OR3_X1    g571(.A1(new_n736_), .A2(G78gat), .A3(new_n666_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n752_), .A2(new_n287_), .A3(new_n753_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G78gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT110), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n731_), .A2(new_n497_), .A3(new_n734_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n695_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n443_), .A2(new_n514_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT111), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n675_), .A2(new_n783_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n514_), .B1(new_n788_), .B2(new_n443_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT112), .ZN(G1336gat));
  INV_X1    g590(.A(new_n788_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G92gat), .B1(new_n792_), .B2(new_n452_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n684_), .A2(new_n515_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n784_), .B2(new_n794_), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n695_), .A2(new_n357_), .A3(new_n783_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G99gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n792_), .A2(new_n523_), .A3(new_n357_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n797_), .A2(new_n798_), .B1(KEYINPUT113), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(KEYINPUT113), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n695_), .A2(new_n287_), .A3(new_n783_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(G106gat), .A3(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n792_), .A2(new_n524_), .A3(new_n287_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT114), .ZN(new_n809_));
  INV_X1    g608(.A(new_n806_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n803_), .A2(G106gat), .A3(new_n810_), .A4(new_n804_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n807_), .A2(new_n814_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1339gat));
  NAND3_X1  g615(.A1(new_n681_), .A2(new_n497_), .A3(new_n631_), .ZN(new_n817_));
  OR3_X1    g616(.A1(new_n817_), .A2(KEYINPUT54), .A3(new_n595_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n817_), .B2(new_n595_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  NAND2_X1  g621(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n576_), .B1(new_n532_), .B2(new_n472_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n578_), .A2(new_n582_), .A3(new_n575_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n822_), .B1(new_n827_), .B2(new_n573_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n584_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n574_), .B1(new_n577_), .B2(new_n583_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n573_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(KEYINPUT117), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n825_), .A2(new_n826_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT55), .A3(new_n573_), .A4(new_n574_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n828_), .A2(new_n830_), .A3(new_n833_), .A4(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n591_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(KEYINPUT56), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n599_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n598_), .A2(new_n604_), .A3(new_n601_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n630_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n625_), .A2(new_n626_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n625_), .A2(new_n626_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT119), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n732_), .A2(new_n847_), .A3(new_n842_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n838_), .A2(new_n839_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(new_n837_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n836_), .A2(KEYINPUT56), .A3(new_n837_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT120), .A3(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n586_), .A2(new_n837_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n849_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(KEYINPUT121), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n857_), .B2(KEYINPUT121), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n681_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT116), .B1(new_n631_), .B2(new_n855_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n734_), .A2(new_n864_), .A3(new_n856_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n827_), .A2(new_n822_), .A3(new_n573_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n831_), .B2(new_n832_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n830_), .A2(new_n835_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n591_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT118), .B1(new_n871_), .B2(KEYINPUT56), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n850_), .A2(new_n873_), .A3(new_n851_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n866_), .B1(new_n875_), .B2(new_n853_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n592_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n566_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n873_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n880_));
  AOI211_X1 g679(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n836_), .C2(new_n837_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n853_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n863_), .A2(new_n865_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n877_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n879_), .B1(new_n884_), .B2(new_n637_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n878_), .A2(new_n885_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n821_), .B(new_n498_), .C1(new_n862_), .C2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n857_), .A2(KEYINPUT121), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT58), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n571_), .A3(new_n859_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n885_), .A3(new_n878_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n821_), .B1(new_n892_), .B2(new_n498_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n820_), .B1(new_n888_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n452_), .A2(new_n443_), .A3(new_n686_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n498_), .B1(new_n862_), .B2(new_n886_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n820_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT59), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n897_), .A2(G113gat), .A3(new_n734_), .A4(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n334_), .B1(new_n900_), .B2(new_n631_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1340gat));
  NAND3_X1  g703(.A1(new_n897_), .A2(new_n595_), .A3(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G120gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n899_), .A2(new_n896_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n330_), .B1(new_n731_), .B2(KEYINPUT60), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n330_), .A2(KEYINPUT60), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n907_), .A2(KEYINPUT123), .A3(new_n908_), .A4(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n906_), .A2(new_n914_), .ZN(G1341gat));
  NAND4_X1  g714(.A1(new_n897_), .A2(G127gat), .A3(new_n497_), .A4(new_n901_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n331_), .B1(new_n900_), .B2(new_n498_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1342gat));
  NAND4_X1  g717(.A1(new_n897_), .A2(G134gat), .A3(new_n571_), .A4(new_n901_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n332_), .B1(new_n900_), .B2(new_n566_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1343gat));
  AOI21_X1  g720(.A(new_n685_), .B1(new_n898_), .B2(new_n820_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n452_), .A2(new_n443_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n631_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n611_), .ZN(G1344gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n731_), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g727(.A1(new_n924_), .A2(new_n498_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT61), .B(G155gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  NOR3_X1   g730(.A1(new_n924_), .A2(new_n559_), .A3(new_n681_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n922_), .A2(new_n637_), .A3(new_n923_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n559_), .B2(new_n933_), .ZN(G1347gat));
  XOR2_X1   g733(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n820_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n898_), .A2(KEYINPUT122), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n887_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n684_), .A2(new_n431_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n686_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n939_), .A2(new_n631_), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(G169gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n936_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n403_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n894_), .A2(new_n734_), .A3(new_n942_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(G169gat), .A3(new_n935_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n946_), .A2(new_n947_), .A3(new_n949_), .ZN(G1348gat));
  NOR2_X1   g749(.A1(new_n939_), .A2(new_n943_), .ZN(new_n951_));
  AOI21_X1  g750(.A(G176gat), .B1(new_n951_), .B2(new_n595_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n941_), .A2(new_n660_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n899_), .A2(new_n666_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n954_), .A2(new_n322_), .A3(new_n731_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n952_), .B1(new_n953_), .B2(new_n955_), .ZN(G1349gat));
  NOR2_X1   g755(.A1(new_n954_), .A2(new_n498_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n317_), .B1(new_n957_), .B2(new_n953_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n498_), .A2(new_n391_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n958_), .B1(new_n951_), .B2(new_n959_), .ZN(G1350gat));
  NAND3_X1  g759(.A1(new_n951_), .A2(new_n637_), .A3(new_n290_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n939_), .A2(new_n681_), .A3(new_n943_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n311_), .B2(new_n962_), .ZN(G1351gat));
  NAND2_X1  g762(.A1(new_n922_), .A2(new_n940_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n631_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n965_), .A2(KEYINPUT125), .A3(new_n208_), .ZN(new_n966_));
  XOR2_X1   g765(.A(KEYINPUT125), .B(G197gat), .Z(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n965_), .B2(new_n967_), .ZN(G1352gat));
  AOI211_X1 g767(.A(new_n685_), .B(new_n941_), .C1(new_n898_), .C2(new_n820_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n595_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g770(.A(KEYINPUT63), .B(G211gat), .C1(new_n969_), .C2(new_n497_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n964_), .A2(new_n498_), .ZN(new_n973_));
  XOR2_X1   g772(.A(KEYINPUT63), .B(G211gat), .Z(new_n974_));
  AOI21_X1  g773(.A(new_n972_), .B1(new_n973_), .B2(new_n974_), .ZN(G1354gat));
  INV_X1    g774(.A(G218gat), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n969_), .A2(new_n976_), .A3(new_n637_), .ZN(new_n977_));
  INV_X1    g776(.A(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n976_), .B1(new_n969_), .B2(new_n571_), .ZN(new_n979_));
  OAI21_X1  g778(.A(KEYINPUT126), .B1(new_n978_), .B2(new_n979_), .ZN(new_n980_));
  INV_X1    g779(.A(new_n979_), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n981_), .A2(new_n982_), .A3(new_n977_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n980_), .A2(new_n983_), .ZN(G1355gat));
endmodule


