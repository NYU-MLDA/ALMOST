//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT66), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  AND2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n204_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n209_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n205_), .A2(KEYINPUT66), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT67), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n212_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT9), .ZN(new_n222_));
  AND2_X1   g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n222_), .B1(KEYINPUT9), .B2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G106gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232_));
  NOR4_X1   g031(.A1(new_n227_), .A2(new_n228_), .A3(new_n232_), .A4(G106gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n226_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n219_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n210_), .A2(new_n211_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n238_), .A2(new_n239_), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(G99gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n241_), .A3(new_n230_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n225_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  OR2_X1    g044(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n246_), .A2(new_n237_), .B1(new_n241_), .B2(new_n230_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n242_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n212_), .A2(new_n218_), .A3(new_n249_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT8), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n235_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n254_));
  INV_X1    g053(.A(G57gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G64gat), .ZN(new_n256_));
  INV_X1    g055(.A(G64gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(G57gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n254_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G71gat), .B(G78gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(G57gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n255_), .A2(G64gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT11), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n260_), .A2(KEYINPUT11), .A3(new_n262_), .A4(new_n263_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n253_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n253_), .A2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n203_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n252_), .A2(new_n245_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n235_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n265_), .A2(new_n267_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n266_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT71), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(new_n284_), .A3(KEYINPUT12), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n253_), .B2(new_n270_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n203_), .B1(new_n253_), .B2(new_n270_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n273_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G120gat), .B(G148gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G176gat), .B(G204gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n290_), .B(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT13), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(KEYINPUT13), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT73), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT34), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G29gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G43gat), .B(G50gat), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n305_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n276_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT15), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n307_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT15), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n253_), .A2(new_n314_), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT35), .B(new_n303_), .C1(new_n309_), .C2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n309_), .A2(new_n315_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n303_), .B(KEYINPUT35), .Z(new_n319_));
  AOI22_X1  g118(.A1(new_n316_), .A2(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT36), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G190gat), .B(G218gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT75), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G134gat), .B(G162gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n303_), .A2(KEYINPUT35), .ZN(new_n327_));
  INV_X1    g126(.A(new_n314_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n276_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n253_), .A2(new_n311_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n327_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT74), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n320_), .A2(new_n321_), .A3(new_n326_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n321_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(KEYINPUT36), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n329_), .A2(new_n330_), .A3(new_n319_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n331_), .B2(KEYINPUT74), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n334_), .B(new_n335_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n333_), .A2(new_n339_), .A3(KEYINPUT37), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT37), .B1(new_n333_), .B2(new_n339_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G127gat), .B(G155gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT16), .ZN(new_n345_));
  XOR2_X1   g144(.A(G183gat), .B(G211gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT76), .B(G8gat), .ZN(new_n348_));
  INV_X1    g147(.A(G1gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT14), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G22gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G8gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G231gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n284_), .ZN(new_n359_));
  AOI211_X1 g158(.A(new_n343_), .B(new_n347_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n358_), .B(new_n270_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n347_), .B(KEYINPUT17), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n342_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n301_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT96), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  OR2_X1    g170(.A1(G197gat), .A2(G204gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(KEYINPUT21), .A3(new_n373_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n377_), .A2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT84), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(KEYINPUT23), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT92), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT92), .B1(new_n394_), .B2(new_n390_), .ZN(new_n395_));
  INV_X1    g194(.A(G169gat), .ZN(new_n396_));
  INV_X1    g195(.A(G176gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G169gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(new_n397_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n384_), .B2(KEYINPUT23), .ZN(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT26), .B(G190gat), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT25), .B(G183gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT24), .B1(new_n396_), .B2(new_n397_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G169gat), .A2(G176gat), .ZN(new_n409_));
  MUX2_X1   g208(.A(new_n408_), .B(KEYINPUT24), .S(new_n409_), .Z(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n382_), .B1(new_n401_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(G183gat), .ZN(new_n413_));
  INV_X1    g212(.A(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n403_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(G176gat), .B1(KEYINPUT85), .B2(KEYINPUT22), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G169gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT26), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n404_), .B2(KEYINPUT83), .ZN(new_n422_));
  INV_X1    g221(.A(G183gat), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n423_), .A2(KEYINPUT82), .A3(KEYINPUT25), .ZN(new_n424_));
  OR3_X1    g223(.A1(new_n423_), .A2(KEYINPUT81), .A3(KEYINPUT82), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT25), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(KEYINPUT81), .B2(new_n423_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n422_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n388_), .A3(new_n410_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n419_), .A2(new_n430_), .A3(new_n382_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT20), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n371_), .B1(new_n412_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n419_), .A2(new_n430_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n381_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n371_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n401_), .A2(new_n382_), .A3(new_n411_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT18), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G64gat), .B(G92gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n369_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n433_), .A2(new_n439_), .A3(KEYINPUT96), .A4(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n412_), .A2(new_n432_), .A3(new_n371_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n444_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT27), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n440_), .A2(new_n444_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n446_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n453_), .A2(KEYINPUT27), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT90), .ZN(new_n457_));
  OR3_X1    g256(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G141gat), .A2(G148gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT89), .A3(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n465_), .B2(KEYINPUT89), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n461_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n465_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n462_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n458_), .A2(new_n459_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT1), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n460_), .B(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n457_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n474_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(new_n470_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n485_), .A3(KEYINPUT90), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT29), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G22gat), .B(G50gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT28), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n489_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n382_), .B1(G228gat), .B2(G233gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n469_), .A2(new_n471_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n498_), .A2(new_n483_), .B1(new_n481_), .B2(new_n474_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n381_), .B1(new_n499_), .B2(new_n488_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G228gat), .A3(G233gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n492_), .B1(new_n493_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n502_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n497_), .A2(new_n495_), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n504_), .A2(new_n492_), .A3(new_n493_), .A4(new_n505_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n456_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G1gat), .B(G29gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(G57gat), .B(G85gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND2_X1  g314(.A1(G225gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G127gat), .B(G134gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G120gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n499_), .A2(KEYINPUT93), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n482_), .A2(new_n485_), .A3(new_n519_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n519_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n480_), .A2(new_n486_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT4), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n516_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n516_), .A3(new_n526_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n524_), .A2(KEYINPUT95), .A3(new_n516_), .A4(new_n526_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n515_), .B1(new_n531_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n516_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n529_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n530_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n515_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G99gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n435_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G227gat), .A2(G233gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT86), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT30), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n552_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT87), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT87), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n557_), .A3(new_n554_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n519_), .B(KEYINPUT31), .Z(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(KEYINPUT87), .A3(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n545_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n510_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n543_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n453_), .A2(new_n454_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n534_), .A2(new_n535_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n568_), .A2(KEYINPUT33), .A3(new_n542_), .A4(new_n541_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n516_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n570_), .B(new_n515_), .C1(new_n516_), .C2(new_n527_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n448_), .A2(new_n449_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n446_), .A2(KEYINPUT32), .ZN(new_n574_));
  MUX2_X1   g373(.A(new_n573_), .B(new_n440_), .S(new_n574_), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n544_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n509_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n509_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n456_), .A2(new_n545_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n560_), .A2(new_n562_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n564_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n356_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G229gat), .A2(G233gat), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n311_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n355_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n308_), .A3(new_n353_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n356_), .A2(KEYINPUT77), .A3(new_n308_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n587_), .B1(new_n593_), .B2(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT80), .ZN(new_n595_));
  XOR2_X1   g394(.A(G113gat), .B(G141gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(G169gat), .B(G197gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n594_), .A2(KEYINPUT80), .A3(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n583_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n368_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n349_), .A3(new_n544_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n333_), .A2(new_n339_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n583_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n604_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n300_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n365_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n545_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT97), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n608_), .A2(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(new_n456_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n606_), .A2(new_n619_), .A3(new_n348_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT98), .ZN(new_n621_));
  OAI21_X1  g420(.A(G8gat), .B1(new_n615_), .B2(new_n456_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT39), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n615_), .B2(new_n582_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT99), .Z(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT41), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT41), .ZN(new_n629_));
  INV_X1    g428(.A(new_n606_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n630_), .A2(G15gat), .A3(new_n582_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n628_), .A2(new_n629_), .A3(KEYINPUT100), .A4(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1326gat));
  OAI21_X1  g435(.A(G22gat), .B1(new_n615_), .B2(new_n509_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n509_), .A2(G22gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n639_), .B1(new_n630_), .B2(new_n640_), .ZN(G1327gat));
  NAND2_X1  g440(.A1(new_n610_), .A2(new_n365_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT106), .ZN(new_n643_));
  INV_X1    g442(.A(new_n300_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n605_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n544_), .ZN(new_n647_));
  XOR2_X1   g446(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n648_));
  INV_X1    g447(.A(new_n342_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n582_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n651_), .B2(new_n564_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(KEYINPUT43), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n579_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n507_), .A2(new_n537_), .A3(new_n543_), .A4(new_n508_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n455_), .B2(new_n452_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n582_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n650_), .A2(new_n456_), .A3(new_n545_), .A4(new_n509_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n342_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n655_), .B1(new_n661_), .B2(KEYINPUT102), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n654_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n613_), .A2(new_n366_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT103), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666_));
  INV_X1    g465(.A(new_n664_), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n666_), .B(new_n667_), .C1(new_n654_), .C2(new_n662_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n648_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT43), .B1(new_n652_), .B2(new_n653_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n661_), .A2(KEYINPUT102), .A3(new_n655_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT44), .B(new_n664_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n663_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n664_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n669_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n544_), .A2(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n647_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(new_n646_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n680_), .A2(G36gat), .A3(new_n456_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n681_), .B(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n669_), .A2(new_n676_), .A3(new_n619_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n669_), .A2(new_n676_), .A3(KEYINPUT107), .A4(new_n619_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G36gat), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT46), .B(new_n684_), .C1(new_n688_), .C2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n681_), .B(new_n682_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n689_), .A2(G36gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(new_n687_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(G1329gat));
  NAND3_X1  g495(.A1(new_n677_), .A2(G43gat), .A3(new_n650_), .ZN(new_n697_));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n680_), .B2(new_n582_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1330gat));
  AOI21_X1  g503(.A(G50gat), .B1(new_n646_), .B2(new_n579_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n579_), .A2(G50gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n677_), .B2(new_n706_), .ZN(G1331gat));
  NOR2_X1   g506(.A1(new_n583_), .A2(new_n612_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n708_), .A2(new_n366_), .A3(new_n644_), .A4(new_n342_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n255_), .B1(new_n709_), .B2(new_n545_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT110), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n611_), .A2(new_n366_), .A3(new_n604_), .A4(new_n301_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT111), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n545_), .A2(new_n255_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n713_), .B2(new_n714_), .ZN(G1332gat));
  AOI21_X1  g514(.A(new_n257_), .B1(new_n713_), .B2(new_n619_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n619_), .A2(new_n257_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n709_), .B2(new_n718_), .ZN(G1333gat));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n650_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(G71gat), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G71gat), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n582_), .A2(G71gat), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n722_), .A2(new_n723_), .B1(new_n709_), .B2(new_n724_), .ZN(G1334gat));
  NAND2_X1  g524(.A1(new_n713_), .A2(new_n579_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G78gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT50), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n509_), .A2(G78gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n709_), .B2(new_n729_), .ZN(G1335gat));
  INV_X1    g529(.A(new_n301_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n643_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n708_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n220_), .A3(new_n544_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n663_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n644_), .A2(new_n365_), .A3(new_n604_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n736_), .A2(new_n545_), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n738_), .B2(new_n220_), .ZN(G1336gat));
  NAND3_X1  g538(.A1(new_n734_), .A2(new_n221_), .A3(new_n619_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n736_), .A2(new_n456_), .A3(new_n737_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n221_), .ZN(G1337gat));
  NOR2_X1   g541(.A1(new_n736_), .A2(new_n737_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n241_), .B1(new_n743_), .B2(new_n650_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT113), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n650_), .A2(new_n229_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT114), .B1(new_n734_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  AOI21_X1  g552(.A(new_n230_), .B1(new_n743_), .B2(new_n579_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n734_), .A2(new_n230_), .A3(new_n579_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  AND4_X1   g561(.A1(new_n366_), .A2(new_n300_), .A3(new_n342_), .A4(new_n604_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT54), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT122), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n285_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n253_), .A2(new_n270_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n285_), .A2(new_n287_), .A3(new_n767_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n766_), .A2(KEYINPUT55), .B1(new_n768_), .B2(new_n203_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n289_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n289_), .A2(KEYINPUT117), .A3(new_n770_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n769_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n295_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n587_), .B(new_n600_), .C1(new_n593_), .C2(new_n585_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n585_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n593_), .B2(new_n585_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n780_), .B1(new_n782_), .B2(new_n600_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT119), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n273_), .A2(new_n289_), .A3(new_n296_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n780_), .B(new_n786_), .C1(new_n782_), .C2(new_n600_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n784_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n784_), .A2(KEYINPUT120), .A3(new_n785_), .A4(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n295_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT121), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n295_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n779_), .B(new_n792_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n765_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n342_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n779_), .A2(new_n792_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n795_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT121), .A3(new_n793_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n800_), .A2(new_n802_), .A3(KEYINPUT122), .A4(KEYINPUT58), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(new_n799_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n784_), .A2(new_n787_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n297_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n602_), .A2(new_n785_), .A3(new_n603_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n811_));
  INV_X1    g610(.A(new_n776_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n776_), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n807_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n805_), .B1(new_n815_), .B2(new_n610_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n810_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n811_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n814_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n807_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n610_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT57), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n804_), .A2(new_n816_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n764_), .B1(new_n365_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n510_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n582_), .A2(new_n545_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n612_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT59), .B1(new_n824_), .B2(new_n828_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n804_), .A2(new_n816_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n804_), .A2(new_n816_), .A3(KEYINPUT124), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n822_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n764_), .B1(new_n839_), .B2(new_n365_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n829_), .A2(KEYINPUT123), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n829_), .A2(KEYINPUT123), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n834_), .B(KEYINPUT125), .C1(new_n840_), .C2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n822_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n366_), .B1(new_n849_), .B2(new_n838_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n844_), .B1(new_n850_), .B2(new_n764_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT125), .B1(new_n851_), .B2(new_n834_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n847_), .A2(new_n852_), .A3(new_n604_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n833_), .B1(new_n853_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n300_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n831_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n851_), .A2(new_n301_), .A3(new_n834_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n859_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n831_), .A2(new_n861_), .A3(new_n366_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n847_), .A2(new_n852_), .A3(new_n365_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1342gat));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n831_), .A2(new_n865_), .A3(new_n610_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n847_), .A2(new_n852_), .A3(new_n342_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n650_), .A2(new_n545_), .A3(new_n509_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n825_), .A2(new_n456_), .A3(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n604_), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n871_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n731_), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g673(.A1(new_n870_), .A2(new_n365_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n870_), .B2(new_n342_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n609_), .A2(G162gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n870_), .B2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n563_), .A2(new_n456_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n509_), .B(new_n881_), .C1(new_n850_), .C2(new_n764_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882_), .B2(new_n604_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n884_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n882_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n399_), .A3(new_n612_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(new_n886_), .A3(new_n888_), .ZN(G1348gat));
  AOI21_X1  g688(.A(G176gat), .B1(new_n887_), .B2(new_n644_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n824_), .A2(new_n579_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n881_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n731_), .A2(new_n397_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n891_), .B2(new_n893_), .ZN(G1349gat));
  NOR3_X1   g693(.A1(new_n882_), .A2(new_n406_), .A3(new_n365_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n366_), .A3(new_n881_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n413_), .B2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n882_), .B2(new_n342_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n610_), .A2(new_n405_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n882_), .B2(new_n899_), .ZN(G1351gat));
  NOR4_X1   g699(.A1(new_n824_), .A2(new_n657_), .A3(new_n456_), .A4(new_n650_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n612_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n301_), .ZN(new_n904_));
  INV_X1    g703(.A(G204gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(KEYINPUT126), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n904_), .B(new_n906_), .ZN(G1353gat));
  AOI21_X1  g706(.A(new_n365_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT127), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n901_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n910_), .B(new_n911_), .Z(G1354gat));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n901_), .A2(new_n913_), .A3(new_n610_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n901_), .A2(new_n649_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n913_), .ZN(G1355gat));
endmodule


