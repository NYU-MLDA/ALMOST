//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n206_));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n212_), .A2(KEYINPUT65), .A3(G85gat), .A4(G92gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT10), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT10), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n211_), .A2(new_n216_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n224_), .A3(new_n223_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT6), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n232_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT8), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n222_), .A2(new_n231_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n220_), .A3(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .A3(new_n232_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n210_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT12), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n208_), .A2(new_n209_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n211_), .A2(new_n216_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n235_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n257_), .B2(new_n220_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n226_), .A2(G99gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n224_), .A2(KEYINPUT10), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT64), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n262_));
  AOI21_X1  g061(.A(G106gat), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n264_));
  OAI22_X1  g063(.A1(KEYINPUT8), .A2(new_n258_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n234_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT66), .B1(new_n234_), .B2(new_n235_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n269_), .B2(new_n220_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n253_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT67), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G230gat), .A2(G233gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n244_), .A2(new_n249_), .A3(new_n210_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n252_), .A2(new_n273_), .A3(new_n274_), .A4(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n275_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G148gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G176gat), .B(G204gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(G120gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n276_), .A2(new_n279_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT70), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n285_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n287_), .A2(new_n289_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(KEYINPUT13), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT71), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G141gat), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G197gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT77), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G29gat), .B(G36gat), .Z(new_n313_));
  INV_X1    g112(.A(G43gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G29gat), .B(G36gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G43gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(G50gat), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n317_), .ZN(new_n319_));
  INV_X1    g118(.A(G50gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G1gat), .B(G8gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT74), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G15gat), .B(G22gat), .ZN(new_n324_));
  INV_X1    g123(.A(G1gat), .ZN(new_n325_));
  INV_X1    g124(.A(G8gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT14), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n323_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n322_), .A2(KEYINPUT74), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n322_), .A2(KEYINPUT74), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n318_), .B(new_n321_), .C1(new_n329_), .C2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n323_), .A2(new_n328_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n315_), .A2(G50gat), .A3(new_n317_), .ZN(new_n337_));
  AOI21_X1  g136(.A(G50gat), .B1(new_n315_), .B2(new_n317_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n335_), .B(new_n336_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(KEYINPUT75), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT75), .B1(new_n334_), .B2(new_n339_), .ZN(new_n342_));
  OAI211_X1 g141(.A(KEYINPUT76), .B(new_n312_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n329_), .A2(new_n333_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n321_), .A2(new_n318_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT15), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n321_), .A2(KEYINPUT15), .A3(new_n318_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n351_), .B2(new_n345_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n344_), .B1(new_n352_), .B2(new_n311_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n334_), .A2(new_n339_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n311_), .B1(new_n356_), .B2(new_n340_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n310_), .B(new_n343_), .C1(new_n353_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n345_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n311_), .A3(new_n334_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT76), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n312_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n310_), .B1(new_n364_), .B2(new_n343_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n359_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n303_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370_));
  INV_X1    g169(.A(G113gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G113gat), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n372_), .A2(G120gat), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(G120gat), .B1(new_n372_), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  OR2_X1    g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT82), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT1), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n380_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n378_), .B(new_n379_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n381_), .B(KEYINPUT83), .C1(G155gat), .C2(G162gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n379_), .A2(KEYINPUT3), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n378_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n379_), .A2(KEYINPUT3), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n392_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n377_), .B1(new_n389_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT95), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT95), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n404_), .A3(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n389_), .A2(new_n399_), .A3(new_n377_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n400_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT94), .B1(new_n408_), .B2(KEYINPUT4), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n410_));
  NOR4_X1   g209(.A1(new_n407_), .A2(new_n400_), .A3(new_n410_), .A4(new_n401_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n369_), .B(new_n406_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n368_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G1gat), .B(G29gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT99), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n412_), .A2(new_n413_), .A3(new_n419_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G204gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(G197gat), .ZN(new_n426_));
  OR2_X1    g225(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(G197gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT21), .B1(new_n307_), .B2(new_n425_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n429_), .B2(new_n307_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G211gat), .B(G218gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(G197gat), .B1(new_n427_), .B2(new_n428_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT85), .B1(new_n438_), .B2(new_n433_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n432_), .A2(new_n436_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT21), .B1(new_n437_), .B2(new_n441_), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n442_), .A2(new_n430_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT25), .B(G183gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT26), .B(G190gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT78), .ZN(new_n449_));
  NOR3_X1   g248(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G176gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n305_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G183gat), .ZN(new_n457_));
  INV_X1    g256(.A(G190gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT23), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT23), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(G183gat), .A3(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n446_), .A2(new_n447_), .A3(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n449_), .A2(new_n456_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(G176gat), .B1(new_n466_), .B2(KEYINPUT22), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT22), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n454_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n459_), .A2(new_n471_), .A3(new_n461_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n460_), .A2(KEYINPUT80), .A3(G183gat), .A4(G190gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n457_), .A2(new_n458_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n470_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n465_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n445_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n445_), .A2(new_n478_), .A3(KEYINPUT92), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n472_), .A2(new_n473_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n448_), .A3(new_n456_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT89), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n485_), .A2(new_n488_), .A3(new_n448_), .A4(new_n456_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n462_), .A2(KEYINPUT91), .A3(new_n475_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT91), .B1(new_n462_), .B2(new_n475_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT22), .B(G169gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT90), .B1(new_n493_), .B2(new_n453_), .ZN(new_n494_));
  MUX2_X1   g293(.A(KEYINPUT90), .B(new_n494_), .S(new_n455_), .Z(new_n495_));
  AOI22_X1  g294(.A1(new_n487_), .A2(new_n489_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n445_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n484_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT19), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n483_), .A2(KEYINPUT93), .A3(new_n498_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n445_), .A2(new_n478_), .A3(KEYINPUT92), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT92), .B1(new_n445_), .B2(new_n478_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n501_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n496_), .A2(new_n497_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT20), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n440_), .A2(new_n444_), .A3(new_n477_), .A4(new_n465_), .ZN(new_n510_));
  OAI211_X1 g309(.A(KEYINPUT20), .B(new_n510_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n500_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT18), .B(G64gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G92gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G8gat), .B(G36gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT32), .ZN(new_n517_));
  AND4_X1   g316(.A1(new_n502_), .A2(new_n509_), .A3(new_n512_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT98), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n511_), .A2(new_n500_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n455_), .A2(KEYINPUT90), .ZN(new_n521_));
  OAI221_X1 g320(.A(new_n521_), .B1(new_n454_), .B2(new_n494_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n486_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT20), .B1(new_n523_), .B2(new_n445_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT97), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT97), .B(KEYINPUT20), .C1(new_n523_), .C2(new_n445_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n483_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n520_), .B1(new_n528_), .B2(new_n500_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n519_), .B1(new_n529_), .B2(new_n517_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n517_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n525_), .A2(new_n524_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n501_), .B1(new_n532_), .B2(new_n527_), .ZN(new_n533_));
  OAI211_X1 g332(.A(KEYINPUT98), .B(new_n531_), .C1(new_n533_), .C2(new_n520_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n518_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n414_), .A2(KEYINPUT99), .A3(new_n420_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n424_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n483_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n538_), .A2(new_n503_), .B1(new_n500_), .B2(new_n511_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n516_), .B1(new_n539_), .B2(new_n502_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n509_), .A2(new_n502_), .A3(new_n512_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n516_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n368_), .B(new_n406_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n408_), .A2(new_n369_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n420_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT33), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n423_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n412_), .A2(KEYINPUT33), .A3(new_n413_), .A4(new_n419_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n544_), .A2(new_n547_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n537_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G228gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n389_), .B2(new_n399_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n556_), .B2(new_n497_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n556_), .A2(new_n497_), .A3(new_n554_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G78gat), .B(G106gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT88), .B1(new_n558_), .B2(new_n559_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n389_), .A2(new_n555_), .A3(new_n399_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G22gat), .B(G50gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT28), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n564_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n389_), .A2(new_n399_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n553_), .B(new_n445_), .C1(new_n572_), .C2(new_n555_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n561_), .B1(new_n573_), .B2(new_n557_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n574_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n562_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n565_), .A2(new_n570_), .A3(new_n564_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n563_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n561_), .A4(new_n560_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G15gat), .B(G43gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G99gat), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n465_), .A2(new_n477_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n465_), .B2(new_n477_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G227gat), .A2(G233gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT30), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT81), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT31), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT31), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n596_), .A3(new_n600_), .A4(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n377_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n377_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n552_), .A2(new_n580_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT27), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n542_), .B1(new_n533_), .B2(new_n520_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(KEYINPUT27), .C1(new_n541_), .C2(new_n542_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n424_), .A2(new_n536_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n580_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n604_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n614_), .A2(new_n602_), .B1(new_n579_), .B2(new_n576_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n611_), .B(new_n612_), .C1(new_n613_), .C2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n606_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT34), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(KEYINPUT35), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n349_), .A2(new_n350_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT72), .ZN(new_n623_));
  OAI211_X1 g422(.A(KEYINPUT35), .B(new_n620_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n244_), .A2(new_n249_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n346_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n627_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n621_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT73), .B(G190gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(G218gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n636_), .B1(new_n630_), .B2(new_n637_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n618_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n630_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n635_), .A3(new_n634_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT37), .A3(new_n638_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n253_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(new_n345_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G183gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(G211gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n650_), .B(new_n651_), .Z(new_n652_));
  INV_X1    g451(.A(KEYINPUT17), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n648_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n654_), .B2(new_n648_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n645_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n617_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n367_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n612_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(KEYINPUT100), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n424_), .A2(KEYINPUT100), .A3(new_n536_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n661_), .A2(G1gat), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT102), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n366_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n298_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n639_), .A2(new_n640_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n658_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n617_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n662_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G1gat), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n669_), .A2(new_n670_), .A3(new_n683_), .A4(KEYINPUT38), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n673_), .A2(new_n674_), .A3(new_n682_), .A4(new_n684_), .ZN(G1324gat));
  INV_X1    g484(.A(new_n661_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n608_), .A2(new_n610_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n326_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT39), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n680_), .A2(new_n687_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G8gat), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT39), .B(new_n326_), .C1(new_n680_), .C2(new_n687_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n605_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n680_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT41), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n686_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n580_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n680_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT42), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1327gat));
  NOR3_X1   g505(.A1(new_n639_), .A2(new_n640_), .A3(new_n657_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n617_), .A2(new_n677_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G29gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n662_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n676_), .A2(new_n657_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n617_), .B2(new_n645_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n645_), .ZN(new_n716_));
  AOI211_X1 g515(.A(KEYINPUT43), .B(new_n716_), .C1(new_n606_), .C2(new_n616_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n712_), .B(new_n713_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n712_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n702_), .B1(new_n537_), .B2(new_n551_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n614_), .A2(new_n579_), .A3(new_n576_), .A4(new_n602_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n580_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n687_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n605_), .A2(new_n720_), .B1(new_n723_), .B2(new_n612_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n724_), .B2(new_n716_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n617_), .A2(new_n714_), .A3(new_n645_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n718_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n665_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n711_), .B1(new_n730_), .B2(G29gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT104), .B(new_n709_), .C1(new_n729_), .C2(new_n665_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n710_), .B1(new_n731_), .B2(new_n732_), .ZN(G1328gat));
  INV_X1    g532(.A(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n708_), .A2(new_n734_), .A3(new_n687_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT45), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n729_), .A2(new_n687_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT105), .B1(new_n737_), .B2(G36gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n739_), .B(new_n734_), .C1(new_n729_), .C2(new_n687_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT46), .B(new_n736_), .C1(new_n738_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  AOI21_X1  g544(.A(new_n314_), .B1(new_n729_), .B2(new_n696_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n708_), .A2(new_n314_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n696_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g548(.A1(new_n708_), .A2(new_n320_), .A3(new_n702_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n729_), .A2(new_n702_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n320_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n724_), .A2(new_n675_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n303_), .A3(new_n679_), .ZN(new_n754_));
  INV_X1    g553(.A(G57gat), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n612_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(KEYINPUT107), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n724_), .B2(new_n675_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n659_), .A2(new_n299_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT106), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT108), .Z(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n665_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n756_), .B1(new_n765_), .B2(new_n755_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n767_), .A3(new_n687_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G64gat), .B1(new_n754_), .B2(new_n611_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT48), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n772_), .A3(new_n696_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G71gat), .B1(new_n754_), .B2(new_n605_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1334gat));
  INV_X1    g575(.A(G78gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n764_), .A2(new_n777_), .A3(new_n702_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G78gat), .B1(new_n754_), .B2(new_n580_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT50), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1335gat));
  NAND2_X1  g580(.A1(new_n303_), .A2(new_n707_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n665_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n725_), .A2(new_n726_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n298_), .A2(new_n657_), .A3(new_n675_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(G85gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n784_), .B1(new_n788_), .B2(new_n662_), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n783_), .B2(new_n687_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n787_), .A2(new_n687_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G92gat), .ZN(G1337gat));
  OAI211_X1 g591(.A(new_n783_), .B(new_n696_), .C1(new_n230_), .C2(new_n229_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n787_), .A2(new_n696_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT109), .B(new_n793_), .C1(new_n794_), .C2(new_n224_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n702_), .A3(new_n786_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n785_), .A2(KEYINPUT111), .A3(new_n702_), .A4(new_n786_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(G106gat), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n783_), .A2(new_n223_), .A3(new_n702_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT110), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n783_), .A2(new_n806_), .A3(new_n223_), .A4(new_n702_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n799_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n800_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n803_), .A2(new_n808_), .A3(new_n812_), .A4(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  NAND3_X1  g613(.A1(new_n659_), .A2(new_n366_), .A3(new_n298_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT54), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n276_), .A2(KEYINPUT112), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n276_), .B2(KEYINPUT112), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n252_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n821_), .A2(new_n278_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n819_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT113), .B(KEYINPUT56), .C1(new_n823_), .C2(new_n285_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n286_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n365_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n358_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n276_), .A2(KEYINPUT112), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT55), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n821_), .A2(new_n278_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n276_), .A2(KEYINPUT112), .A3(new_n818_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n285_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n824_), .B(new_n827_), .C1(KEYINPUT56), .C2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n312_), .B1(new_n356_), .B2(new_n340_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n309_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n311_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT114), .A3(new_n308_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n352_), .A2(new_n312_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n364_), .A2(new_n309_), .A3(new_n343_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n292_), .A2(new_n294_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n678_), .B1(new_n836_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n817_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n844_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n291_), .A2(new_n850_), .A3(new_n293_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n286_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT113), .B1(new_n823_), .B2(new_n285_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n855_), .B2(new_n824_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT115), .B(KEYINPUT57), .C1(new_n856_), .C2(new_n678_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n849_), .A2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n285_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n833_), .A2(new_n854_), .A3(new_n834_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n286_), .A3(new_n845_), .A4(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n833_), .A2(new_n834_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n825_), .B1(new_n864_), .B2(KEYINPUT56), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT58), .A3(new_n845_), .A4(new_n860_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n645_), .A3(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n858_), .A2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n816_), .B1(new_n868_), .B2(new_n657_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n615_), .B(new_n611_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT118), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n870_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n872_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n867_), .A2(KEYINPUT116), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n863_), .A2(new_n645_), .A3(new_n866_), .A4(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n858_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n858_), .A2(new_n878_), .A3(KEYINPUT117), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n658_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n874_), .B1(new_n883_), .B2(new_n816_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n675_), .B(new_n873_), .C1(new_n884_), .C2(new_n870_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n371_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n884_), .A2(KEYINPUT119), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n888_), .B(new_n874_), .C1(new_n883_), .C2(new_n816_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n675_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n371_), .B2(new_n890_), .ZN(G1340gat));
  OR2_X1    g690(.A1(new_n884_), .A2(new_n870_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n303_), .A3(new_n873_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G120gat), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895_));
  AOI21_X1  g694(.A(G120gat), .B1(new_n299_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT120), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n895_), .B2(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT121), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n901_), .B(new_n898_), .C1(new_n887_), .C2(new_n889_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n894_), .A2(new_n900_), .A3(new_n902_), .ZN(G1341gat));
  INV_X1    g702(.A(G127gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n657_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n905_));
  OAI211_X1 g704(.A(G127gat), .B(new_n873_), .C1(new_n884_), .C2(new_n870_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n904_), .A2(new_n905_), .B1(new_n907_), .B2(new_n657_), .ZN(G1342gat));
  AND2_X1   g707(.A1(new_n892_), .A2(new_n873_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n645_), .A2(G134gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT122), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n678_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n912_));
  INV_X1    g711(.A(G134gat), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n909_), .A2(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1343gat));
  AOI21_X1  g713(.A(new_n721_), .B1(new_n883_), .B2(new_n816_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n666_), .A2(new_n687_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n675_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(G141gat), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n918_), .B(new_n920_), .ZN(G1344gat));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n303_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT124), .B(G148gat), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n922_), .B(new_n924_), .ZN(G1345gat));
  NAND2_X1  g724(.A1(new_n917_), .A2(new_n657_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT61), .B(G155gat), .Z(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT125), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n926_), .B(new_n928_), .ZN(G1346gat));
  AOI21_X1  g728(.A(G162gat), .B1(new_n917_), .B2(new_n678_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n645_), .A2(G162gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n917_), .B2(new_n931_), .ZN(G1347gat));
  AND4_X1   g731(.A1(new_n615_), .A2(new_n869_), .A3(new_n687_), .A4(new_n666_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n305_), .B1(new_n933_), .B2(new_n675_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n934_), .A2(KEYINPUT62), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(new_n493_), .A3(new_n675_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(KEYINPUT62), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(G1348gat));
  AOI21_X1  g737(.A(G176gat), .B1(new_n933_), .B2(new_n299_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n702_), .B1(new_n883_), .B2(new_n816_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n665_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n941_), .A2(G176gat), .A3(new_n303_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n939_), .B1(new_n940_), .B2(new_n942_), .ZN(G1349gat));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n657_), .A3(new_n941_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n940_), .A2(KEYINPUT126), .A3(new_n657_), .A4(new_n941_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n946_), .A2(new_n457_), .A3(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n446_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n933_), .A2(new_n657_), .A3(new_n949_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n948_), .A2(new_n950_), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n933_), .A2(new_n678_), .A3(new_n447_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n933_), .A2(new_n645_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n458_), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n662_), .A2(new_n611_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n858_), .A2(new_n878_), .A3(KEYINPUT117), .ZN(new_n956_));
  AOI21_X1  g755(.A(KEYINPUT117), .B1(new_n858_), .B2(new_n878_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n956_), .A2(new_n957_), .A3(new_n657_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n816_), .ZN(new_n959_));
  OAI211_X1 g758(.A(new_n613_), .B(new_n955_), .C1(new_n958_), .C2(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(KEYINPUT127), .B1(new_n915_), .B2(new_n955_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n675_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(G197gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n960_), .A2(new_n961_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n915_), .A2(KEYINPUT127), .A3(new_n955_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n968_), .A2(new_n307_), .A3(new_n675_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n965_), .A2(new_n969_), .ZN(G1352gat));
  NAND3_X1  g769(.A1(new_n968_), .A2(new_n429_), .A3(new_n303_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n303_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n972_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n971_), .B1(new_n425_), .B2(new_n973_), .ZN(G1353gat));
  OR2_X1    g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n975_), .B1(new_n968_), .B2(new_n657_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(KEYINPUT63), .B(G211gat), .ZN(new_n977_));
  AOI211_X1 g776(.A(new_n658_), .B(new_n977_), .C1(new_n966_), .C2(new_n967_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n976_), .A2(new_n978_), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n968_), .B2(new_n678_), .ZN(new_n980_));
  INV_X1    g779(.A(G218gat), .ZN(new_n981_));
  AOI211_X1 g780(.A(new_n981_), .B(new_n716_), .C1(new_n966_), .C2(new_n967_), .ZN(new_n982_));
  NOR2_X1   g781(.A1(new_n980_), .A2(new_n982_), .ZN(G1355gat));
endmodule


