//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT85), .B1(G183gat), .B2(G190gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT23), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT85), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n202_), .B(new_n205_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT83), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT83), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n220_), .A2(KEYINPUT84), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n207_), .B(new_n222_), .C1(new_n220_), .C2(KEYINPUT84), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n210_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT94), .B(G204gat), .Z(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(G197gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT93), .B(G197gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(G204gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT21), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n225_), .A2(G197gat), .B1(new_n227_), .B2(G204gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT21), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n231_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n234_), .B1(new_n230_), .B2(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n224_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n207_), .B1(G183gat), .B2(G190gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n202_), .B(KEYINPUT97), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n203_), .B(KEYINPUT98), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n238_), .B(new_n239_), .C1(new_n241_), .C2(G176gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n213_), .B(KEYINPUT96), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(new_n218_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n212_), .A3(new_n222_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n242_), .B1(new_n208_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT20), .B1(new_n246_), .B2(new_n236_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT19), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n237_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n224_), .A2(new_n236_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT20), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n246_), .B2(new_n236_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G64gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(G92gat), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT103), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(KEYINPUT103), .A3(new_n260_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT27), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n249_), .B1(new_n237_), .B2(new_n247_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n252_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n260_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(new_n264_), .A3(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n269_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n261_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n265_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G225gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT100), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n278_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n278_), .B2(KEYINPUT2), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT89), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT90), .Z(new_n283_));
  NOR2_X1   g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT3), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT87), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n284_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n288_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(KEYINPUT1), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n291_), .B(new_n292_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT99), .ZN(new_n301_));
  INV_X1    g100(.A(new_n299_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n290_), .A2(new_n302_), .A3(new_n295_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n296_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(KEYINPUT99), .A3(new_n302_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(KEYINPUT4), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n277_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n275_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT0), .ZN(new_n315_));
  INV_X1    g114(.A(G57gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G85gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n313_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n271_), .A2(new_n274_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n296_), .A2(KEYINPUT29), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(new_n325_), .B2(new_n236_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n236_), .A3(new_n324_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G78gat), .B(G106gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT95), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n328_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n329_), .B1(new_n334_), .B2(new_n326_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n296_), .A2(KEYINPUT29), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n296_), .B2(KEYINPUT29), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G22gat), .B(G50gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n341_), .A3(new_n339_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n344_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n333_), .B(new_n336_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n335_), .A2(new_n331_), .A3(new_n345_), .A4(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n224_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT86), .ZN(new_n354_));
  XOR2_X1   g153(.A(G71gat), .B(G99gat), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  NOR2_X1   g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n224_), .B(KEYINPUT30), .ZN(new_n358_));
  INV_X1    g157(.A(new_n356_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n299_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G15gat), .B(G43gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT31), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n352_), .A2(new_n356_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n302_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n361_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n350_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n348_), .B(new_n349_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n323_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n311_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n277_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n373_), .A2(new_n320_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n273_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n378_));
  NOR4_X1   g177(.A1(new_n310_), .A2(KEYINPUT33), .A3(new_n312_), .A4(new_n319_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT101), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n376_), .B(KEYINPUT101), .C1(new_n378_), .C2(new_n379_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n256_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n385_), .A2(KEYINPUT102), .ZN(new_n386_));
  INV_X1    g185(.A(new_n384_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n385_), .A2(KEYINPUT102), .B1(new_n387_), .B2(new_n268_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n321_), .A2(new_n322_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(new_n383_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n350_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n369_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n372_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G183gat), .B(G211gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G127gat), .B(G155gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT17), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT77), .B(G22gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G15gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n405_));
  XOR2_X1   g204(.A(KEYINPUT78), .B(G1gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT79), .B(G8gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G1gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G8gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n409_), .A2(new_n410_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n404_), .A2(new_n408_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G1gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(G8gat), .B1(new_n417_), .B2(new_n411_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G231gat), .A2(G233gat), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n415_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n413_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(G8gat), .A3(new_n411_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n421_), .A2(new_n422_), .B1(G231gat), .B2(G233gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G57gat), .B(G64gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT11), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427_));
  AND2_X1   g226(.A1(KEYINPUT69), .A2(G71gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(KEYINPUT69), .A2(G71gat), .ZN(new_n429_));
  INV_X1    g228(.A(G78gat), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G64gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G57gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n316_), .A2(G64gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT11), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n427_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT69), .A2(G71gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT69), .A2(G71gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(G78gat), .A3(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(new_n437_), .C1(KEYINPUT11), .C2(new_n425_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(KEYINPUT70), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n426_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(KEYINPUT70), .ZN(new_n445_));
  INV_X1    g244(.A(new_n435_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(new_n427_), .A3(new_n437_), .A4(new_n441_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n426_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n402_), .B1(new_n424_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n451_), .B2(new_n424_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n444_), .A2(KEYINPUT72), .A3(new_n449_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT72), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n445_), .A2(new_n448_), .A3(new_n447_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n448_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n424_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT17), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n401_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n454_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT81), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n459_), .A2(new_n466_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n453_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G232gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT34), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT35), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G29gat), .B(G36gat), .Z(new_n475_));
  XOR2_X1   g274(.A(G43gat), .B(G50gat), .Z(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT15), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT65), .B1(new_n485_), .B2(new_n480_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT64), .B(G92gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n318_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT10), .B(G99gat), .Z(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n488_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  XOR2_X1   g297(.A(G85gat), .B(G92gat), .Z(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT66), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT66), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT67), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n508_));
  NOR4_X1   g307(.A1(new_n508_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n504_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n498_), .B(new_n499_), .C1(new_n510_), .C2(new_n487_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n485_), .A2(new_n480_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n504_), .B(new_n512_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n498_), .B1(new_n513_), .B2(new_n499_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n514_), .B2(KEYINPUT68), .ZN(new_n515_));
  INV_X1    g314(.A(new_n499_), .ZN(new_n516_));
  INV_X1    g315(.A(G99gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n506_), .A2(new_n517_), .A3(new_n495_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n508_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n505_), .A2(KEYINPUT67), .A3(new_n506_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n519_), .A2(new_n520_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n516_), .B1(new_n521_), .B2(new_n512_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n498_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n497_), .B1(new_n515_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n479_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI22_X1  g326(.A1(new_n525_), .A2(new_n477_), .B1(KEYINPUT35), .B2(new_n471_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n474_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n497_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n499_), .A2(new_n498_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n488_), .B2(new_n521_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n513_), .A2(new_n499_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT8), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n534_), .B2(new_n523_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n477_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n537_), .A2(new_n538_), .B1(new_n473_), .B2(new_n472_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n474_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n526_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n529_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G134gat), .B(G162gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT75), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n215_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G218gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT36), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n548_), .A2(KEYINPUT76), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n529_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n548_), .B2(KEYINPUT76), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n396_), .A2(new_n469_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n537_), .B2(new_n450_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n462_), .A2(KEYINPUT12), .A3(new_n525_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n523_), .B1(new_n522_), .B2(new_n498_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n536_), .A3(new_n511_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n450_), .A3(new_n497_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .A4(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n525_), .A2(new_n451_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(KEYINPUT71), .A3(new_n562_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n450_), .B1(new_n561_), .B2(new_n497_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n558_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G120gat), .B(G148gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(G204gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT5), .B(G176gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n563_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n573_), .B(KEYINPUT73), .Z(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n575_), .A2(new_n577_), .A3(KEYINPUT74), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n563_), .A2(new_n569_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n576_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n582_), .B2(new_n574_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n555_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT74), .B1(new_n575_), .B2(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n579_), .A3(new_n574_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n586_), .A3(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G169gat), .ZN(new_n590_));
  INV_X1    g389(.A(G197gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n415_), .A2(new_n418_), .A3(new_n478_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n477_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G229gat), .A2(G233gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n594_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n538_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n421_), .A2(new_n422_), .A3(new_n477_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n593_), .B1(new_n598_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n600_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n597_), .B1(new_n603_), .B2(new_n595_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n479_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n596_), .A3(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n606_), .A3(new_n592_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n602_), .A2(KEYINPUT82), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT82), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n593_), .C1(new_n598_), .C2(new_n601_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n588_), .A2(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT105), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT105), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n554_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n390_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n548_), .A2(KEYINPUT37), .A3(new_n551_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n468_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n612_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n396_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n406_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n390_), .A3(new_n627_), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n628_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n618_), .A2(new_n629_), .A3(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n407_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n271_), .A2(new_n274_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n624_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n554_), .A2(new_n634_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(G8gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(G8gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n369_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n624_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n615_), .A2(new_n643_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(new_n645_), .B2(G15gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n624_), .A2(new_n649_), .A3(new_n350_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G22gat), .B1(new_n616_), .B2(new_n393_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT42), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(KEYINPUT42), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n396_), .A2(new_n623_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n553_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n468_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n390_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n613_), .A2(new_n469_), .A3(new_n614_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n620_), .A2(new_n621_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n396_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n380_), .A2(new_n381_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n394_), .B1(new_n665_), .B2(new_n383_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n664_), .B(new_n661_), .C1(new_n666_), .C2(new_n372_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n660_), .B1(new_n663_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT44), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n669_), .A2(G29gat), .A3(new_n390_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n659_), .B1(new_n670_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n633_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n658_), .A2(new_n675_), .A3(new_n634_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(KEYINPUT46), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  INV_X1    g482(.A(new_n680_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n679_), .B(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n685_), .B2(new_n677_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n682_), .A2(new_n686_), .ZN(G1329gat));
  NAND3_X1  g486(.A1(new_n655_), .A2(new_n643_), .A3(new_n657_), .ZN(new_n688_));
  INV_X1    g487(.A(G43gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT108), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n669_), .A2(G43gat), .A3(new_n643_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n672_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT47), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n691_), .B(new_n695_), .C1(new_n672_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n658_), .B2(new_n350_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n669_), .A2(G50gat), .A3(new_n350_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n673_), .ZN(G1331gat));
  AND3_X1   g499(.A1(new_n554_), .A2(new_n588_), .A3(new_n611_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n617_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n611_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n396_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(new_n611_), .C1(new_n666_), .C2(new_n372_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n705_), .A2(new_n588_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n622_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n390_), .A2(new_n316_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n703_), .B1(new_n710_), .B2(new_n711_), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n432_), .B1(new_n701_), .B2(new_n634_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT48), .Z(new_n714_));
  INV_X1    g513(.A(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n432_), .A3(new_n634_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n701_), .B2(new_n643_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n718_), .A3(new_n643_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  AOI21_X1  g521(.A(new_n430_), .B1(new_n701_), .B2(new_n350_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n715_), .A2(new_n430_), .A3(new_n350_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1335gat));
  NAND2_X1  g526(.A1(new_n663_), .A2(new_n667_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n588_), .A2(new_n469_), .A3(new_n611_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT111), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n728_), .A2(KEYINPUT112), .A3(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n318_), .B1(new_n735_), .B2(new_n390_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n705_), .A2(new_n707_), .A3(new_n588_), .A4(new_n657_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n737_), .A2(G85gat), .A3(new_n617_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1336gat));
  INV_X1    g538(.A(new_n737_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G92gat), .B1(new_n740_), .B2(new_n634_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n633_), .A2(new_n490_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n735_), .B2(new_n742_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n494_), .A3(new_n643_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n369_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n517_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT51), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n744_), .B(new_n748_), .C1(new_n745_), .C2(new_n517_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1338gat));
  NAND2_X1  g549(.A1(new_n350_), .A2(new_n495_), .ZN(new_n751_));
  OR3_X1    g550(.A1(new_n737_), .A2(KEYINPUT113), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n737_), .B2(new_n751_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n495_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n731_), .B2(new_n393_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI221_X1 g557(.A(new_n755_), .B1(KEYINPUT114), .B2(KEYINPUT52), .C1(new_n731_), .C2(new_n393_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n754_), .A2(new_n758_), .A3(new_n762_), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  NAND3_X1  g563(.A1(new_n584_), .A2(new_n587_), .A3(new_n611_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT115), .B1(new_n622_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n622_), .A2(new_n765_), .A3(KEYINPUT115), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n622_), .A2(new_n765_), .A3(KEYINPUT115), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT54), .B1(new_n771_), .B2(new_n766_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n599_), .A2(KEYINPUT117), .A3(new_n605_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n597_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n599_), .A2(new_n600_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n592_), .B1(new_n778_), .B2(new_n596_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n607_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(new_n574_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n559_), .A2(new_n562_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n558_), .A2(KEYINPUT116), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n783_), .A2(KEYINPUT55), .A3(new_n557_), .A4(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n563_), .A2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n557_), .A2(KEYINPUT55), .A3(new_n559_), .A4(new_n562_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n784_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n581_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n581_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n782_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n782_), .B(KEYINPUT58), .C1(new_n793_), .C2(new_n792_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n661_), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n781_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT118), .B(new_n781_), .C1(new_n578_), .C2(new_n583_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n608_), .A2(new_n574_), .A3(new_n610_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n801_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n656_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n798_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n656_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n469_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n773_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n634_), .A2(new_n617_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n371_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n811_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n806_), .B(new_n798_), .C1(new_n808_), .C2(new_n816_), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n805_), .C2(new_n656_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n469_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n773_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n814_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n821_), .B2(new_n811_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n611_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(new_n824_), .A3(new_n704_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(new_n588_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n820_), .B(new_n814_), .C1(KEYINPUT60), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n588_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G120gat), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(KEYINPUT60), .B2(new_n829_), .ZN(G1341gat));
  OAI21_X1  g631(.A(G127gat), .B1(new_n822_), .B2(new_n469_), .ZN(new_n833_));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n821_), .A2(new_n834_), .A3(new_n468_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1342gat));
  OAI21_X1  g635(.A(G134gat), .B1(new_n822_), .B2(new_n662_), .ZN(new_n837_));
  INV_X1    g636(.A(G134gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n821_), .A2(new_n838_), .A3(new_n553_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1343gat));
  OAI21_X1  g639(.A(new_n769_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n771_), .A2(KEYINPUT54), .A3(new_n766_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n808_), .A2(new_n816_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n808_), .A2(new_n816_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n798_), .A2(new_n806_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n843_), .B1(new_n847_), .B2(new_n469_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n848_), .A2(new_n370_), .A3(new_n813_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n704_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n588_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT120), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NAND2_X1  g653(.A1(new_n849_), .A2(new_n468_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  AOI21_X1  g656(.A(G162gat), .B1(new_n849_), .B2(new_n553_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n661_), .A2(G162gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT121), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n849_), .B2(new_n860_), .ZN(G1347gat));
  NAND3_X1  g660(.A1(new_n634_), .A2(new_n617_), .A3(new_n643_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT122), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n350_), .B(new_n863_), .C1(new_n773_), .C2(new_n809_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n704_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G169gat), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n868_), .B(new_n869_), .C1(new_n241_), .C2(new_n865_), .ZN(G1348gat));
  AOI21_X1  g669(.A(G176gat), .B1(new_n864_), .B2(new_n588_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n848_), .A2(new_n350_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n863_), .A2(new_n204_), .A3(new_n827_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  INV_X1    g673(.A(new_n863_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n872_), .A2(new_n468_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G183gat), .B1(new_n876_), .B2(new_n877_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n469_), .A2(new_n243_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n878_), .A2(new_n879_), .B1(new_n864_), .B2(new_n880_), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n864_), .A2(new_n553_), .A3(new_n218_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n864_), .A2(new_n661_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n215_), .ZN(G1351gat));
  NOR3_X1   g683(.A1(new_n370_), .A2(new_n633_), .A3(new_n390_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT124), .B1(new_n820_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  INV_X1    g686(.A(new_n885_), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n887_), .B(new_n888_), .C1(new_n819_), .C2(new_n773_), .ZN(new_n889_));
  OAI211_X1 g688(.A(G197gat), .B(new_n704_), .C1(new_n886_), .C2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n887_), .B1(new_n848_), .B2(new_n888_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n820_), .A2(KEYINPUT124), .A3(new_n885_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(G197gat), .A4(new_n704_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n704_), .B1(new_n886_), .B2(new_n889_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n591_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n891_), .A2(new_n896_), .A3(new_n898_), .ZN(G1352gat));
  AOI21_X1  g698(.A(G204gat), .B1(new_n894_), .B2(new_n588_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n827_), .B(new_n225_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1353gat));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT126), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n469_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n894_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n894_), .B2(new_n905_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1354gat));
  NAND2_X1  g707(.A1(new_n894_), .A2(new_n553_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT127), .B(G218gat), .Z(new_n910_));
  NOR2_X1   g709(.A1(new_n662_), .A2(new_n910_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n909_), .A2(new_n910_), .B1(new_n894_), .B2(new_n911_), .ZN(G1355gat));
endmodule


