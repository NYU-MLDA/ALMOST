//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_;
  INV_X1    g000(.A(KEYINPUT109), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT2), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G141gat), .A3(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT88), .ZN(new_n207_));
  AOI22_X1  g006(.A1(new_n204_), .A2(new_n206_), .B1(new_n207_), .B2(KEYINPUT3), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n209_), .B(new_n210_), .C1(new_n207_), .C2(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n212_), .B(KEYINPUT88), .C1(G141gat), .C2(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT89), .B1(new_n208_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  INV_X1    g015(.A(G155gat), .ZN(new_n217_));
  INV_X1    g016(.A(G162gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n208_), .A2(KEYINPUT89), .A3(new_n214_), .ZN(new_n224_));
  OR2_X1    g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(KEYINPUT1), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n219_), .A2(new_n228_), .A3(new_n220_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n225_), .A3(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G141gat), .B(G148gat), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n226_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  INV_X1    g033(.A(G134gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT85), .B(G127gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n226_), .A3(new_n232_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT4), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n233_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT105), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n240_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT106), .B(KEYINPUT0), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G1gat), .B(G29gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT108), .ZN(new_n257_));
  INV_X1    g056(.A(new_n255_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n258_), .A3(new_n249_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT108), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n250_), .A2(new_n260_), .A3(new_n255_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT19), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT23), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(G183gat), .A3(G190gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n268_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT100), .B(KEYINPUT24), .Z(new_n273_));
  OR2_X1    g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n271_), .B(new_n272_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT101), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n276_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT25), .B(G183gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT99), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G190gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .A4(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT22), .B(G169gat), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n278_), .B(KEYINPUT102), .Z(new_n289_));
  NAND3_X1  g088(.A1(new_n267_), .A2(new_n269_), .A3(KEYINPUT83), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT83), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n266_), .A2(new_n291_), .A3(KEYINPUT23), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n288_), .B(new_n289_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n285_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n298_));
  INV_X1    g097(.A(G204gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT92), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n299_), .A2(G197gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n298_), .A2(KEYINPUT92), .A3(new_n299_), .A4(new_n300_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT21), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT94), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G211gat), .A2(G218gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT94), .B1(new_n313_), .B2(new_n308_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(G204gat), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n299_), .A2(G197gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n318_), .A2(new_n320_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(KEYINPUT93), .A3(new_n319_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n307_), .A2(new_n315_), .A3(new_n323_), .A4(new_n325_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n312_), .A2(new_n314_), .A3(KEYINPUT95), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT95), .B1(new_n312_), .B2(new_n314_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n324_), .A2(new_n319_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n297_), .A2(new_n332_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n306_), .A2(KEYINPUT21), .B1(new_n314_), .B2(new_n312_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n321_), .B(KEYINPUT93), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n334_), .A2(new_n335_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n274_), .A2(KEYINPUT24), .A3(new_n278_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n274_), .A2(KEYINPUT24), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(new_n339_), .B2(G190gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n281_), .B(new_n340_), .C1(new_n283_), .C2(KEYINPUT82), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n293_), .A2(new_n337_), .A3(new_n338_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n271_), .A2(new_n272_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n278_), .B(new_n288_), .C1(new_n343_), .C2(new_n295_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT20), .B1(new_n336_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n265_), .B1(new_n333_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n297_), .A2(new_n332_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n336_), .A2(new_n346_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n349_), .A2(KEYINPUT20), .A3(new_n264_), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n353_));
  XOR2_X1   g152(.A(KEYINPUT104), .B(G8gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT103), .B(KEYINPUT18), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n333_), .A2(new_n347_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(new_n265_), .ZN(new_n363_));
  AND4_X1   g162(.A1(KEYINPUT20), .A2(new_n349_), .A3(new_n265_), .A4(new_n350_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT32), .B(new_n361_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n262_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n352_), .B(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n259_), .A2(KEYINPUT107), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT33), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n242_), .A2(new_n245_), .A3(new_n244_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n240_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n255_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT33), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n259_), .A2(KEYINPUT107), .A3(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n367_), .A2(new_n369_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n366_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n377_), .B(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n226_), .B2(new_n232_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n385_), .A2(new_n336_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n224_), .A2(new_n225_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n389_), .A2(new_n215_), .A3(new_n222_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n232_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT29), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n386_), .B1(new_n392_), .B2(new_n332_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n383_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n387_), .B1(new_n385_), .B2(new_n336_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n386_), .A3(new_n332_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n382_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n381_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT96), .B1(new_n388_), .B2(new_n393_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT96), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n383_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT97), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n381_), .A2(new_n397_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n399_), .A2(new_n401_), .A3(KEYINPUT97), .A4(new_n383_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT98), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n404_), .A2(KEYINPUT98), .A3(new_n405_), .A4(new_n406_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n398_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n342_), .A2(new_n344_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n345_), .A2(KEYINPUT30), .ZN(new_n418_));
  INV_X1    g217(.A(new_n413_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n342_), .A2(new_n344_), .A3(new_n414_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G43gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n417_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n412_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n415_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n419_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n422_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n412_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n417_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n426_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n238_), .B(KEYINPUT31), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n426_), .A2(new_n432_), .A3(new_n433_), .A4(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n376_), .A2(new_n411_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n409_), .A2(new_n410_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n398_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n439_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n411_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n367_), .A2(KEYINPUT27), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n359_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n352_), .A2(new_n361_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(KEYINPUT27), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(new_n262_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n440_), .B1(new_n447_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G15gat), .B(G22gat), .ZN(new_n455_));
  INV_X1    g254(.A(G1gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G1gat), .B(G8gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G29gat), .B(G36gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n461_), .B(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n461_), .A2(new_n464_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n464_), .B(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n468_), .B2(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470_));
  MUX2_X1   g269(.A(new_n465_), .B(new_n469_), .S(new_n470_), .Z(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT80), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT78), .B(KEYINPUT79), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G169gat), .B(G197gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n471_), .A2(new_n477_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n202_), .B1(new_n454_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G190gat), .B(G218gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G134gat), .B(G162gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT36), .ZN(new_n489_));
  INV_X1    g288(.A(G85gat), .ZN(new_n490_));
  INV_X1    g289(.A(G92gat), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT9), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT6), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT9), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G85gat), .B(G92gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT10), .B(G99gat), .ZN(new_n500_));
  OAI221_X1 g299(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .C1(G106gat), .C2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n496_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT65), .ZN(new_n503_));
  AND2_X1   g302(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n504_));
  NOR2_X1   g303(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  MUX2_X1   g306(.A(new_n506_), .B(new_n504_), .S(new_n507_), .Z(new_n508_));
  AOI21_X1  g307(.A(new_n499_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AOI211_X1 g310(.A(KEYINPUT8), .B(new_n499_), .C1(new_n508_), .C2(new_n502_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n501_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(new_n464_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n468_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n518_), .A2(new_n519_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n488_), .A2(KEYINPUT36), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n514_), .A2(new_n526_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n489_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT37), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n528_), .B2(KEYINPUT73), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n533_), .B(new_n489_), .C1(new_n529_), .C2(new_n530_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G231gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n461_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G71gat), .B(G78gat), .ZN(new_n543_));
  OR3_X1    g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n543_), .A3(KEYINPUT11), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n539_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT76), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n547_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n537_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  INV_X1    g362(.A(new_n546_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n513_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT12), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n513_), .A2(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n565_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n565_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT68), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT5), .B(G176gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n576_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n573_), .A2(new_n576_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT67), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n581_), .B(KEYINPUT69), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n573_), .A2(KEYINPUT67), .A3(new_n576_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n563_), .B1(new_n584_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n563_), .A3(new_n590_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n562_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n445_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n595_));
  AOI211_X1 g394(.A(new_n398_), .B(new_n439_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n453_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n376_), .A2(new_n411_), .A3(new_n439_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT109), .A3(new_n482_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n484_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n456_), .A3(new_n262_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n602_), .A2(KEYINPUT110), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n454_), .A2(new_n531_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n593_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n591_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n483_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n605_), .A2(new_n561_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n456_), .B1(new_n609_), .B2(new_n262_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n602_), .B1(new_n610_), .B2(new_n603_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT110), .B1(new_n602_), .B2(new_n603_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n611_), .A3(new_n612_), .ZN(G1324gat));
  NAND3_X1  g412(.A1(new_n609_), .A2(KEYINPUT111), .A3(new_n452_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n605_), .A2(new_n561_), .A3(new_n452_), .A4(new_n608_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT111), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(G8gat), .A3(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT112), .B(KEYINPUT39), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n614_), .A2(G8gat), .A3(new_n621_), .A4(new_n617_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n601_), .A2(new_n457_), .A3(new_n452_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(KEYINPUT40), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  INV_X1    g428(.A(G15gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n601_), .A2(new_n630_), .A3(new_n445_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT113), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n609_), .B2(new_n445_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n609_), .B2(new_n443_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT42), .Z(new_n638_));
  NAND3_X1  g437(.A1(new_n601_), .A2(new_n636_), .A3(new_n443_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n607_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n531_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n561_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n484_), .A2(new_n641_), .A3(new_n600_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n262_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT114), .B(KEYINPUT43), .C1(new_n454_), .C2(new_n537_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT114), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n537_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n607_), .A2(new_n561_), .A3(new_n483_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n654_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n262_), .A2(G29gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n646_), .B1(new_n659_), .B2(new_n660_), .ZN(G1328gat));
  NAND3_X1  g460(.A1(new_n657_), .A2(new_n452_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n644_), .A2(G36gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT45), .B1(new_n664_), .B2(new_n452_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n666_));
  INV_X1    g465(.A(new_n452_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n644_), .A2(new_n666_), .A3(G36gat), .A4(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n663_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT115), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT46), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT115), .B(new_n673_), .C1(new_n663_), .C2(new_n669_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1329gat));
  NAND3_X1  g474(.A1(new_n657_), .A2(new_n445_), .A3(new_n658_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G43gat), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n644_), .A2(G43gat), .A3(new_n439_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1330gat));
  NAND2_X1  g480(.A1(new_n659_), .A2(new_n443_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT116), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT116), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n659_), .A2(new_n684_), .A3(new_n443_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(G50gat), .A3(new_n685_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n644_), .A2(G50gat), .A3(new_n411_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n641_), .A2(new_n482_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n599_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n562_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G57gat), .B1(new_n691_), .B2(new_n262_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n605_), .A2(new_n561_), .A3(new_n689_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n262_), .A2(G57gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(G1332gat));
  INV_X1    g494(.A(G64gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n693_), .B2(new_n452_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT48), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n691_), .A2(new_n696_), .A3(new_n452_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n693_), .B2(new_n445_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT49), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n691_), .A2(new_n701_), .A3(new_n445_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1334gat));
  INV_X1    g504(.A(G78gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n691_), .A2(new_n706_), .A3(new_n443_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n693_), .A2(new_n443_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G78gat), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT117), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1335gat));
  NOR3_X1   g513(.A1(new_n690_), .A2(new_n561_), .A3(new_n642_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G85gat), .B1(new_n715_), .B2(new_n262_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n653_), .A2(new_n560_), .A3(new_n689_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n262_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n490_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n716_), .B1(new_n718_), .B2(new_n720_), .ZN(G1336gat));
  AOI21_X1  g520(.A(G92gat), .B1(new_n715_), .B2(new_n452_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n667_), .A2(new_n491_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n718_), .B2(new_n723_), .ZN(G1337gat));
  OAI21_X1  g523(.A(G99gat), .B1(new_n717_), .B2(new_n439_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(KEYINPUT118), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT119), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n439_), .A2(new_n500_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n715_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(KEYINPUT118), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n726_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT51), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n726_), .A2(new_n733_), .A3(new_n729_), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1338gat));
  INV_X1    g534(.A(G106gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n715_), .A2(new_n736_), .A3(new_n443_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n653_), .A2(new_n560_), .A3(new_n443_), .A4(new_n689_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G106gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G106gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n568_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n575_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n573_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n746_), .A2(new_n745_), .A3(new_n575_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n588_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n482_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n582_), .B(KEYINPUT70), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n584_), .A2(new_n590_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n465_), .A2(new_n470_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n469_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n477_), .B(new_n759_), .C1(new_n760_), .C2(new_n470_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n478_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n755_), .A2(new_n757_), .B1(new_n758_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n744_), .B1(new_n764_), .B2(new_n531_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n751_), .B2(KEYINPUT56), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n756_), .B1(new_n751_), .B2(KEYINPUT56), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(KEYINPUT58), .A3(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n751_), .A2(KEYINPUT56), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n584_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n772_), .B2(new_n766_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n769_), .A2(new_n773_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n758_), .A2(new_n763_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n757_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n754_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT57), .A3(new_n642_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n765_), .A2(new_n774_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n560_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(KEYINPUT120), .A2(KEYINPUT54), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT120), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n594_), .A2(new_n483_), .A3(new_n781_), .A4(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n560_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n483_), .B(new_n786_), .C1(new_n606_), .C2(new_n591_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n452_), .A2(new_n719_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n411_), .A3(new_n445_), .A4(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT123), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n789_), .B1(new_n779_), .B2(new_n560_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n796_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n798_));
  INV_X1    g597(.A(new_n794_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n792_), .A4(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n793_), .A2(KEYINPUT59), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n483_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n795_), .A2(new_n800_), .A3(new_n801_), .A4(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n793_), .B2(new_n483_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1340gat));
  NAND4_X1  g605(.A1(new_n795_), .A2(new_n800_), .A3(new_n607_), .A4(new_n801_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT124), .B(G120gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT125), .ZN(new_n810_));
  INV_X1    g609(.A(new_n808_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n641_), .B2(KEYINPUT60), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n797_), .A2(new_n792_), .A3(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(KEYINPUT60), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n793_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n814_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n816_), .A2(KEYINPUT125), .A3(new_n812_), .A4(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n809_), .A2(new_n819_), .ZN(G1341gat));
  INV_X1    g619(.A(G127gat), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n560_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n795_), .A2(new_n800_), .A3(new_n801_), .A4(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n821_), .B1(new_n793_), .B2(new_n560_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1342gat));
  NOR2_X1   g624(.A1(new_n537_), .A2(new_n235_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n795_), .A2(new_n800_), .A3(new_n801_), .A4(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n235_), .B1(new_n793_), .B2(new_n642_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1343gat));
  NOR2_X1   g628(.A1(new_n796_), .A2(new_n444_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n792_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n483_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(new_n209_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n641_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n210_), .ZN(G1345gat));
  NOR2_X1   g634(.A1(new_n831_), .A2(new_n560_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT61), .B(G155gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  NOR3_X1   g637(.A1(new_n831_), .A2(new_n218_), .A3(new_n537_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n831_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n531_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n218_), .B2(new_n841_), .ZN(G1347gat));
  NOR2_X1   g641(.A1(new_n796_), .A2(new_n443_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n667_), .A2(new_n262_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n445_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(G169gat), .B1(new_n847_), .B2(new_n483_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n843_), .A2(new_n286_), .A3(new_n482_), .A4(new_n846_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n848_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n852_), .B2(new_n849_), .ZN(G1348gat));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n843_), .B(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n855_), .A2(G176gat), .A3(new_n607_), .A4(new_n846_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n287_), .B1(new_n847_), .B2(new_n641_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1349gat));
  NOR3_X1   g657(.A1(new_n847_), .A2(new_n560_), .A3(new_n282_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n855_), .A2(new_n561_), .A3(new_n846_), .ZN(new_n860_));
  INV_X1    g659(.A(G183gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n847_), .B2(new_n537_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n531_), .A2(new_n283_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n847_), .B2(new_n864_), .ZN(G1351gat));
  NAND2_X1  g664(.A1(new_n830_), .A2(new_n844_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n483_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT127), .B(G197gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1352gat));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n641_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n299_), .ZN(G1353gat));
  NOR2_X1   g670(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n872_));
  AND2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n866_), .A2(new_n560_), .A3(new_n872_), .A4(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n866_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n561_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n876_), .B2(new_n872_), .ZN(G1354gat));
  INV_X1    g676(.A(G218gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n866_), .A2(new_n878_), .A3(new_n537_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n531_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n878_), .B2(new_n880_), .ZN(G1355gat));
endmodule


