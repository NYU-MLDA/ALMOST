//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203_));
  INV_X1    g002(.A(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(G57gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G64gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT68), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n207_), .A3(new_n210_), .A4(KEYINPUT11), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n207_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G71gat), .B(G78gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT11), .B1(new_n205_), .B2(new_n207_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT67), .B1(new_n220_), .B2(new_n217_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n212_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n212_), .B1(new_n221_), .B2(new_n219_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n203_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT9), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT64), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n227_), .A2(new_n228_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT6), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT6), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  INV_X1    g042(.A(G106gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n237_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n236_), .A2(new_n247_), .ZN(new_n248_));
  OR3_X1    g047(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n242_), .A2(new_n249_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n228_), .A2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n248_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G57gat), .B(G64gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n210_), .B1(new_n263_), .B2(KEYINPUT11), .ZN(new_n264_));
  INV_X1    g063(.A(new_n211_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n216_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n220_), .A2(KEYINPUT67), .A3(new_n217_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n212_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT69), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n224_), .A2(new_n262_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n235_), .A2(new_n242_), .A3(new_n237_), .A4(new_n246_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n254_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n260_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n269_), .A2(KEYINPUT69), .A3(new_n270_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT69), .B1(new_n269_), .B2(new_n270_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT70), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n262_), .B1(new_n224_), .B2(new_n271_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n202_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n224_), .A2(new_n271_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n288_), .B2(new_n277_), .ZN(new_n289_));
  AOI211_X1 g088(.A(KEYINPUT70), .B(new_n262_), .C1(new_n224_), .C2(new_n271_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n272_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n286_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT71), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n277_), .A2(KEYINPUT72), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n296_), .B(new_n274_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n282_), .B2(KEYINPUT12), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n272_), .A2(new_n286_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n272_), .A2(KEYINPUT73), .A3(new_n286_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n294_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT5), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n294_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(KEYINPUT13), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT13), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n294_), .B2(new_n307_), .ZN(new_n318_));
  AOI211_X1 g117(.A(new_n306_), .B(new_n312_), .C1(new_n287_), .C2(new_n293_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT74), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G57gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328_));
  INV_X1    g127(.A(G141gat), .ZN(new_n329_));
  INV_X1    g128(.A(G148gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT87), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n333_), .A2(new_n337_), .A3(KEYINPUT87), .A4(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n334_), .A2(new_n336_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n331_), .A2(KEYINPUT3), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT2), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n332_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n331_), .A2(KEYINPUT3), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G127gat), .B(G134gat), .Z(new_n355_));
  XOR2_X1   g154(.A(G113gat), .B(G120gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n343_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT95), .A3(new_n357_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n328_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n359_), .B2(KEYINPUT4), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n327_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n362_), .A2(new_n364_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n366_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n373_), .B(new_n326_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT83), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G169gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n376_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G169gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G183gat), .ZN(new_n383_));
  INV_X1    g182(.A(G190gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT23), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(G183gat), .A3(G190gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(KEYINPUT84), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(KEYINPUT23), .C1(new_n383_), .C2(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n378_), .B(new_n382_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT25), .B(G183gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT26), .B(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(new_n387_), .ZN(new_n397_));
  INV_X1    g196(.A(G176gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n381_), .A2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n399_), .A2(KEYINPUT24), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G169gat), .A2(G176gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(KEYINPUT24), .A3(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n396_), .A2(new_n397_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n393_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT85), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n393_), .A2(new_n406_), .A3(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409_));
  INV_X1    g208(.A(G43gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(G15gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT30), .ZN(new_n416_));
  INV_X1    g215(.A(new_n411_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n405_), .A2(new_n407_), .A3(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT31), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n412_), .A2(new_n418_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT31), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n419_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n358_), .B1(new_n422_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n422_), .A2(new_n358_), .A3(new_n427_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n375_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432_));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT28), .B1(new_n354_), .B2(KEYINPUT29), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT28), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n343_), .A2(new_n353_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G22gat), .B(G50gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n435_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n434_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n435_), .A2(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n439_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n435_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n432_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G197gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G204gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT90), .ZN(new_n450_));
  INV_X1    g249(.A(G204gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G197gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT89), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT21), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n452_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT21), .ZN(new_n456_));
  XOR2_X1   g255(.A(G211gat), .B(G218gat), .Z(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(KEYINPUT21), .A3(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(G228gat), .A2(G233gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n437_), .B2(new_n363_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n461_), .B1(new_n363_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n443_), .A2(new_n447_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n469_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G8gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT18), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G64gat), .B(G92gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n408_), .B2(new_n461_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G226gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n396_), .A2(new_n402_), .A3(new_n400_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n483_), .A2(new_n391_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n483_), .B2(new_n391_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n397_), .B1(G183gat), .B2(G190gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n401_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G169gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n398_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n485_), .A2(new_n486_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n482_), .B1(new_n491_), .B2(new_n462_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n479_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n482_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n485_), .A2(new_n486_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n478_), .B1(new_n498_), .B2(new_n461_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n462_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n477_), .B1(new_n494_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n493_), .A3(new_n476_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n500_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n507_), .A2(new_n482_), .B1(new_n479_), .B2(new_n492_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n476_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n482_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n462_), .B(new_n497_), .C1(new_n483_), .C2(new_n391_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n495_), .B1(new_n479_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n477_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n505_), .A2(new_n506_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n431_), .A2(new_n472_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n369_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT33), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n370_), .A2(new_n517_), .A3(new_n327_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n372_), .A2(KEYINPUT4), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n359_), .A2(KEYINPUT4), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n367_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n326_), .B1(new_n372_), .B2(new_n367_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n516_), .A2(new_n518_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n374_), .A2(new_n517_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n524_), .A2(new_n504_), .A3(new_n502_), .A4(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT32), .B(new_n476_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT32), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n508_), .B1(new_n528_), .B2(new_n477_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n375_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n472_), .A2(new_n375_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n531_), .A2(new_n472_), .B1(new_n514_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n534_));
  INV_X1    g333(.A(new_n430_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n428_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n429_), .A2(KEYINPUT86), .A3(new_n430_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n515_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT82), .ZN(new_n540_));
  XOR2_X1   g339(.A(G29gat), .B(G36gat), .Z(new_n541_));
  XOR2_X1   g340(.A(G43gat), .B(G50gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT15), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545_));
  INV_X1    g344(.A(G1gat), .ZN(new_n546_));
  INV_X1    g345(.A(G8gat), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G8gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n544_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n543_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n553_), .B(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n560_), .A2(new_n564_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n540_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT82), .A3(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n539_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT78), .ZN(new_n575_));
  XOR2_X1   g374(.A(G134gat), .B(G162gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n277_), .B2(new_n553_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n262_), .A2(KEYINPUT76), .A3(new_n543_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT79), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n295_), .A2(new_n544_), .A3(new_n297_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n585_), .A2(KEYINPUT77), .A3(new_n587_), .A4(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT35), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  OAI22_X1  g392(.A1(new_n588_), .A2(KEYINPUT35), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n589_), .A2(new_n593_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n581_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n589_), .A2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n593_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n597_), .A2(new_n580_), .A3(new_n598_), .A4(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n579_), .B1(new_n596_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n596_), .B2(KEYINPUT80), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n603_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n551_), .B(new_n608_), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n288_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT81), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n609_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n609_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n607_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n322_), .A2(new_n573_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n546_), .A3(new_n375_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT98), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n321_), .A2(new_n572_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n631_), .A2(KEYINPUT96), .A3(new_n623_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT96), .B1(new_n631_), .B2(new_n623_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n603_), .B(KEYINPUT97), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n539_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n633_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n375_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n630_), .B(new_n638_), .C1(new_n628_), .C2(new_n627_), .ZN(G1324gat));
  XNOR2_X1  g438(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT101), .Z(new_n641_));
  INV_X1    g440(.A(new_n514_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n632_), .A2(new_n642_), .A3(new_n633_), .A4(new_n635_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G8gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT99), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n646_), .A3(G8gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT39), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n650_), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n625_), .A2(G8gat), .A3(new_n514_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n641_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n641_), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n653_), .B(new_n656_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1325gat));
  INV_X1    g457(.A(new_n538_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G15gat), .B1(new_n636_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT41), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n626_), .A2(new_n414_), .A3(new_n538_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n636_), .B2(new_n472_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n667_));
  AND3_X1   g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n472_), .A2(G22gat), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT104), .Z(new_n671_));
  OAI22_X1  g470(.A1(new_n668_), .A2(new_n669_), .B1(new_n625_), .B2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n539_), .A2(new_n673_), .A3(new_n607_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n539_), .A2(new_n607_), .A3(KEYINPUT105), .A4(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n539_), .A2(new_n607_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT43), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n623_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n631_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n637_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n681_), .A2(new_n603_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n321_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n573_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n637_), .A2(G29gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT106), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n686_), .B1(new_n689_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n683_), .B(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n642_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n514_), .A2(G36gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n573_), .A2(new_n688_), .A3(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n695_), .B1(new_n698_), .B2(new_n704_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n694_), .B(new_n703_), .C1(new_n697_), .C2(G36gat), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  NOR2_X1   g506(.A1(new_n535_), .A2(new_n428_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n410_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n685_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n696_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n410_), .B1(new_n689_), .B2(new_n659_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT47), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n711_), .A2(new_n713_), .A3(new_n717_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1330gat));
  OR3_X1    g518(.A1(new_n689_), .A2(G50gat), .A3(new_n472_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n472_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n696_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(KEYINPUT109), .ZN(new_n723_));
  OAI21_X1  g522(.A(G50gat), .B1(new_n722_), .B2(KEYINPUT109), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(G1331gat));
  INV_X1    g524(.A(new_n322_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n681_), .A2(new_n571_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n635_), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n637_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n539_), .A2(new_n571_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n321_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n624_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n206_), .A3(new_n375_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1332gat));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n204_), .A3(new_n642_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G64gat), .B1(new_n729_), .B2(new_n514_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT111), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n740_));
  AND3_X1   g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n741_), .B2(new_n742_), .ZN(G1333gat));
  OAI21_X1  g542(.A(G71gat), .B1(new_n729_), .B2(new_n659_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n747_), .A3(new_n538_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n729_), .B2(new_n472_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(new_n752_), .A3(new_n721_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1335gat));
  NAND3_X1  g553(.A1(new_n726_), .A2(new_n687_), .A3(new_n731_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n225_), .A3(new_n375_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n321_), .A2(new_n572_), .A3(new_n681_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n680_), .A2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n375_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n760_), .B2(new_n225_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n226_), .A3(new_n642_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n759_), .A2(new_n642_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n226_), .ZN(G1337gat));
  NAND2_X1  g563(.A1(new_n243_), .A2(new_n245_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n755_), .A2(new_n708_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n538_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G99gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n768_), .B(new_n770_), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n680_), .A2(new_n721_), .A3(new_n758_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n680_), .A2(KEYINPUT114), .A3(new_n721_), .A4(new_n758_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G106gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT52), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(new_n773_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .A4(new_n775_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n756_), .A2(new_n244_), .A3(new_n721_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NOR4_X1   g586(.A1(new_n642_), .A2(new_n708_), .A3(new_n637_), .A4(new_n721_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n552_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n563_), .B1(new_n557_), .B2(new_n555_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n567_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT119), .B(new_n791_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n319_), .A2(new_n571_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n272_), .A2(KEYINPUT73), .A3(new_n286_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT73), .B1(new_n272_), .B2(new_n286_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n798_), .B1(new_n801_), .B2(new_n301_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n301_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(KEYINPUT55), .C1(new_n800_), .C2(new_n799_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n292_), .B1(new_n301_), .B2(new_n273_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT116), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n292_), .C1(new_n301_), .C2(new_n273_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n802_), .A2(new_n804_), .A3(new_n806_), .A4(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n312_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n809_), .B2(new_n312_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n797_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT118), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n797_), .B(new_n815_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n796_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n603_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n603_), .A2(KEYINPUT57), .ZN(new_n821_));
  INV_X1    g620(.A(new_n791_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT120), .B1(new_n319_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n315_), .A2(new_n824_), .A3(new_n791_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n809_), .B2(new_n312_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n823_), .B(new_n825_), .C1(new_n810_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n606_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n810_), .A2(new_n826_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n830_), .A2(KEYINPUT58), .A3(new_n823_), .A4(new_n825_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n817_), .A2(new_n821_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n681_), .B1(new_n820_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n321_), .A2(new_n728_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n834_), .B2(new_n607_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n321_), .A2(new_n728_), .A3(new_n836_), .A4(new_n606_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(KEYINPUT54), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT115), .B(new_n839_), .C1(new_n834_), .C2(new_n607_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n788_), .B1(new_n833_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n572_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT59), .B(new_n788_), .C1(new_n833_), .C2(new_n841_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n571_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n849_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n321_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n843_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n322_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n851_), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n843_), .A2(new_n856_), .A3(new_n681_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n623_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n634_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n843_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n606_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT121), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n866_), .B(new_n862_), .C1(new_n863_), .C2(new_n860_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n538_), .A2(new_n472_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n642_), .A2(new_n637_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n869_), .B(new_n870_), .C1(new_n833_), .C2(new_n841_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT122), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n572_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G141gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n329_), .A3(new_n572_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n726_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G148gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(new_n330_), .A3(new_n726_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1345gat));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT123), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n872_), .A2(new_n681_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n872_), .B2(new_n681_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n872_), .A2(new_n886_), .A3(new_n861_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n606_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n886_), .B2(new_n890_), .ZN(G1347gat));
  OR2_X1    g690(.A1(new_n833_), .A2(new_n841_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n514_), .A2(new_n375_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n538_), .A2(new_n472_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895_), .B2(new_n571_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n572_), .A3(new_n489_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n897_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n900_), .A3(new_n901_), .ZN(G1348gat));
  OAI21_X1  g701(.A(G176gat), .B1(new_n895_), .B2(new_n322_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n732_), .A2(new_n398_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n895_), .B2(new_n904_), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n895_), .A2(new_n623_), .ZN(new_n906_));
  MUX2_X1   g705(.A(G183gat), .B(new_n394_), .S(new_n906_), .Z(G1350gat));
  OAI211_X1 g706(.A(new_n607_), .B(new_n894_), .C1(new_n833_), .C2(new_n841_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n908_), .A2(new_n909_), .A3(G190gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n908_), .B2(G190gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n861_), .A2(new_n395_), .ZN(new_n912_));
  OAI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n895_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT125), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  OAI221_X1 g714(.A(new_n915_), .B1(new_n895_), .B2(new_n912_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n892_), .A2(new_n869_), .A3(new_n893_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n571_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n448_), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n322_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n451_), .ZN(G1353gat));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(new_n918_), .B2(new_n623_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  OAI211_X1 g725(.A(KEYINPUT127), .B(new_n923_), .C1(new_n918_), .C2(new_n623_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n833_), .A2(new_n841_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n928_), .A2(new_n472_), .A3(new_n538_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  NAND4_X1  g729(.A1(new_n929_), .A2(new_n681_), .A3(new_n893_), .A4(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n918_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n934_), .A2(KEYINPUT126), .A3(new_n681_), .A4(new_n930_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n926_), .A2(new_n927_), .B1(new_n933_), .B2(new_n935_), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n918_), .B2(new_n606_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n634_), .A2(G218gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n918_), .B2(new_n938_), .ZN(G1355gat));
endmodule


