//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT84), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT84), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n205_), .A2(new_n209_), .A3(new_n211_), .A4(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT22), .B(G169gat), .Z(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n204_), .C1(G176gat), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT85), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT85), .B1(new_n215_), .B2(new_n218_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT30), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT88), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G15gat), .B(G43gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT87), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT86), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n228_), .B(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n225_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n219_), .B(new_n220_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT30), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT88), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT31), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241_));
  INV_X1    g040(.A(G120gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT89), .B(G113gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT31), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n233_), .A2(new_n246_), .A3(new_n238_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n240_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n245_), .B1(new_n240_), .B2(new_n247_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n243_), .B(new_n244_), .Z(new_n250_));
  INV_X1    g049(.A(G155gat), .ZN(new_n251_));
  INV_X1    g050(.A(G162gat), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n251_), .A2(new_n252_), .A3(KEYINPUT1), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT1), .B1(new_n251_), .B2(new_n252_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n253_), .B(new_n254_), .C1(G155gat), .C2(G162gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G141gat), .A2(G148gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n256_), .B(KEYINPUT3), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT90), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n261_), .A2(KEYINPUT2), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(KEYINPUT2), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n258_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n263_), .A2(new_n258_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n262_), .A3(new_n264_), .A4(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G155gat), .B(G162gat), .Z(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT91), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n266_), .A2(KEYINPUT91), .A3(new_n267_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n250_), .B(new_n259_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n259_), .B1(new_n269_), .B2(new_n268_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n245_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(KEYINPUT4), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n276_), .A3(new_n245_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT99), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n270_), .A2(new_n274_), .A3(new_n272_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n273_), .A2(KEYINPUT99), .A3(new_n275_), .A4(new_n277_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G85gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT0), .B(G57gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n280_), .A2(new_n287_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n248_), .A2(new_n249_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n271_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G22gat), .B(G50gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G197gat), .B(G204gat), .Z(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT21), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(KEYINPUT21), .ZN(new_n303_));
  XOR2_X1   g102(.A(G211gat), .B(G218gat), .Z(new_n304_));
  OR3_X1    g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n304_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n307_), .B2(KEYINPUT93), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n310_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G78gat), .B(G106gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT94), .Z(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n312_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(KEYINPUT95), .A3(new_n312_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n300_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n316_), .B(new_n314_), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n299_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT27), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n221_), .A2(new_n222_), .A3(new_n307_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT96), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT96), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n329_), .B(KEYINPUT20), .C1(new_n234_), .C2(new_n307_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n307_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n202_), .A2(new_n208_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n211_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT97), .Z(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n214_), .A3(new_n205_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n335_), .A2(new_n218_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n328_), .B(new_n330_), .C1(new_n331_), .C2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT19), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G64gat), .B(G92gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(new_n218_), .A3(new_n331_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(KEYINPUT20), .C1(new_n223_), .C2(new_n331_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(new_n339_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n340_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n340_), .B2(new_n348_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n325_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT103), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT103), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n325_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n347_), .A2(new_n339_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n345_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(KEYINPUT102), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n325_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n349_), .B1(KEYINPUT102), .B2(new_n358_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n352_), .A2(new_n354_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n292_), .A2(new_n324_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n289_), .A2(new_n290_), .B1(new_n356_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n340_), .A2(new_n348_), .A3(new_n364_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT100), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n340_), .A2(KEYINPUT100), .A3(new_n348_), .A4(new_n364_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT101), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n349_), .A2(new_n350_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n270_), .A2(new_n275_), .A3(new_n272_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n273_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n288_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n290_), .A2(KEYINPUT33), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n290_), .A2(KEYINPUT33), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n374_), .B(new_n377_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n366_), .A2(KEYINPUT101), .A3(new_n369_), .A4(new_n370_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n373_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n291_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n382_), .A2(new_n324_), .B1(new_n362_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n248_), .A2(new_n249_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n363_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G230gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT64), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G85gat), .A2(G92gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT9), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G85gat), .ZN(new_n392_));
  INV_X1    g191(.A(G92gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(new_n389_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n388_), .B(new_n391_), .C1(new_n395_), .C2(new_n390_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G99gat), .A2(G106gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT10), .B(G99gat), .Z(new_n402_));
  INV_X1    g201(.A(G106gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n390_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n391_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT64), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n396_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT8), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT65), .ZN(new_n414_));
  AND3_X1   g213(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n399_), .A2(KEYINPUT65), .A3(new_n400_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n409_), .B1(new_n419_), .B2(new_n395_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n401_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n395_), .A2(new_n409_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n408_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G71gat), .B(G78gat), .ZN(new_n425_));
  INV_X1    g224(.A(G57gat), .ZN(new_n426_));
  INV_X1    g225(.A(G64gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G57gat), .A2(G64gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT11), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT11), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n432_), .A3(new_n429_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n425_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G71gat), .B(G78gat), .Z(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(KEYINPUT11), .B2(new_n430_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n424_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(KEYINPUT67), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n437_), .B(new_n408_), .C1(new_n420_), .C2(new_n423_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(KEYINPUT67), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n424_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n447_));
  AND4_X1   g246(.A1(new_n387_), .A2(new_n443_), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n444_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n387_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT66), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT66), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n452_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT5), .B(G176gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G204gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G120gat), .B(G148gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n454_), .A2(new_n456_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n463_), .A2(new_n464_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT68), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT13), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n466_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(G43gat), .B(G50gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(G29gat), .B(G36gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n474_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT15), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT15), .B1(new_n475_), .B2(new_n476_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(KEYINPUT77), .A2(KEYINPUT78), .ZN(new_n480_));
  NOR2_X1   g279(.A1(KEYINPUT77), .A2(KEYINPUT78), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT76), .B(G8gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT75), .B(G1gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(G15gat), .A2(G22gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G15gat), .A2(G22gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n482_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  OR2_X1    g290(.A1(KEYINPUT76), .A2(G8gat), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT75), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT75), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G1gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(KEYINPUT76), .A2(G8gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT14), .ZN(new_n499_));
  INV_X1    g298(.A(new_n482_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n489_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n490_), .A2(new_n491_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n491_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n482_), .B(new_n489_), .C1(new_n498_), .C2(KEYINPUT14), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n479_), .A2(KEYINPUT81), .A3(new_n503_), .A4(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n503_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n475_), .A2(new_n476_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n477_), .A2(new_n478_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n472_), .B(new_n508_), .C1(new_n513_), .C2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n472_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n510_), .A2(new_n512_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n511_), .B1(new_n507_), .B2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT82), .B(G169gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(G197gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT83), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n516_), .A2(new_n520_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n527_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(KEYINPUT83), .A3(new_n525_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n471_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n424_), .A2(new_n511_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n479_), .A2(new_n424_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT71), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT69), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n541_), .A2(new_n542_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n545_), .A2(KEYINPUT69), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(KEYINPUT69), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n252_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT72), .B(G134gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT74), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n549_), .A2(new_n552_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n557_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT73), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n549_), .B2(new_n552_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n534_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n549_), .A2(new_n552_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n562_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n549_), .A2(new_n552_), .A3(new_n559_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT37), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n571_));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n510_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n437_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n575_), .B1(new_n578_), .B2(KEYINPUT17), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(KEYINPUT17), .B2(new_n575_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n578_), .A2(KEYINPUT80), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n570_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n386_), .A2(new_n533_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT104), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n586_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n587_), .A2(KEYINPUT105), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT105), .B1(new_n587_), .B2(new_n588_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n291_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n485_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n386_), .A2(new_n533_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n567_), .A2(new_n568_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT106), .Z(new_n599_));
  NOR3_X1   g398(.A1(new_n597_), .A2(new_n599_), .A3(new_n583_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n592_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(KEYINPUT38), .A3(new_n593_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n596_), .A2(new_n602_), .A3(new_n603_), .ZN(G1324gat));
  OAI21_X1  g403(.A(G8gat), .B1(new_n601_), .B2(new_n362_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT39), .ZN(new_n606_));
  INV_X1    g405(.A(new_n591_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n362_), .A2(new_n484_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n606_), .B(KEYINPUT40), .C1(new_n607_), .C2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n605_), .B(new_n611_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n589_), .A2(new_n590_), .A3(new_n608_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(new_n385_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G15gat), .B1(new_n601_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT41), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n587_), .A2(new_n588_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n619_), .A2(G15gat), .A3(new_n616_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n618_), .A2(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n324_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n600_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT42), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n622_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n619_), .B2(new_n626_), .ZN(G1327gat));
  NOR2_X1   g426(.A1(new_n598_), .A2(new_n582_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n386_), .A2(new_n533_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n291_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n386_), .A2(new_n570_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT43), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n386_), .A2(new_n634_), .A3(new_n570_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n533_), .A3(new_n583_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n636_), .A2(KEYINPUT44), .A3(new_n533_), .A4(new_n583_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(new_n291_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n631_), .B1(new_n642_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g442(.A(new_n362_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n639_), .A2(new_n644_), .A3(new_n640_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n629_), .A2(G36gat), .A3(new_n362_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT45), .Z(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(new_n648_), .A3(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1329gat));
  NAND4_X1  g452(.A1(new_n639_), .A2(G43gat), .A3(new_n385_), .A4(new_n640_), .ZN(new_n654_));
  INV_X1    g453(.A(G43gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n629_), .B2(new_n616_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g457(.A(G50gat), .B1(new_n630_), .B2(new_n623_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n623_), .A2(G50gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n641_), .B2(new_n660_), .ZN(G1331gat));
  NAND2_X1  g460(.A1(new_n386_), .A2(new_n532_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT107), .Z(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n470_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n584_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n426_), .B1(new_n665_), .B2(new_n592_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT108), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n426_), .C1(new_n665_), .C2(new_n592_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n599_), .A2(new_n583_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n530_), .A2(new_n531_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n470_), .A2(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n670_), .A2(new_n386_), .A3(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT109), .B(G57gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n592_), .A2(new_n674_), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n667_), .A2(new_n669_), .B1(new_n673_), .B2(new_n675_), .ZN(G1332gat));
  AOI21_X1  g475(.A(new_n427_), .B1(new_n673_), .B2(new_n644_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT48), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n644_), .A2(new_n427_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n665_), .B2(new_n679_), .ZN(G1333gat));
  INV_X1    g479(.A(G71gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n673_), .B2(new_n385_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT110), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT49), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n665_), .A2(G71gat), .A3(new_n616_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1334gat));
  INV_X1    g485(.A(G78gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n673_), .B2(new_n623_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT50), .Z(new_n689_));
  NAND2_X1  g488(.A1(new_n623_), .A2(new_n687_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n665_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT111), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1335gat));
  AND3_X1   g492(.A1(new_n386_), .A2(new_n634_), .A3(new_n570_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n634_), .B1(new_n386_), .B2(new_n570_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n583_), .B(new_n672_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(new_n392_), .A3(new_n592_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n664_), .A2(new_n291_), .A3(new_n628_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n392_), .ZN(G1336gat));
  NOR3_X1   g498(.A1(new_n696_), .A2(new_n393_), .A3(new_n362_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n664_), .A2(new_n644_), .A3(new_n628_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n393_), .ZN(G1337gat));
  INV_X1    g501(.A(KEYINPUT112), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n696_), .A2(new_n616_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(G99gat), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n703_), .B(G99gat), .C1(new_n696_), .C2(new_n616_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n664_), .A2(new_n628_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n385_), .A2(new_n402_), .ZN(new_n709_));
  OAI22_X1  g508(.A1(new_n705_), .A2(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT51), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712_));
  OAI221_X1 g511(.A(new_n712_), .B1(new_n708_), .B2(new_n709_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1338gat));
  OAI21_X1  g513(.A(G106gat), .B1(new_n696_), .B2(new_n324_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI211_X1 g516(.A(KEYINPUT113), .B(G106gat), .C1(new_n696_), .C2(new_n324_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(KEYINPUT52), .A3(new_n718_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n664_), .A2(new_n403_), .A3(new_n623_), .A4(new_n628_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n715_), .A2(new_n716_), .A3(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT53), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n719_), .A2(new_n725_), .A3(new_n720_), .A4(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  NAND3_X1  g526(.A1(new_n443_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n451_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n448_), .B1(KEYINPUT55), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n447_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n441_), .B1(new_n424_), .B2(new_n438_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n444_), .A2(new_n445_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(KEYINPUT55), .A3(new_n387_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n460_), .B1(new_n730_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT56), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT115), .B1(new_n738_), .B2(KEYINPUT116), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n671_), .A2(new_n462_), .A3(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT115), .B(new_n460_), .C1(new_n730_), .C2(new_n736_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT56), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT117), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n739_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT55), .B1(new_n734_), .B2(new_n387_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n449_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n735_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n460_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(new_n532_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n742_), .A2(new_n743_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n738_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .A4(new_n462_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n517_), .B(new_n508_), .C1(new_n513_), .C2(new_n515_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n472_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n525_), .A3(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n529_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n745_), .A2(new_n755_), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT57), .A3(new_n598_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n761_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n598_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  INV_X1    g565(.A(new_n737_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n462_), .B1(new_n767_), .B2(new_n738_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n759_), .B1(new_n737_), .B2(KEYINPUT56), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n768_), .A2(new_n766_), .A3(new_n769_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n570_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n764_), .A2(new_n765_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n761_), .A2(new_n598_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT118), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n777_), .B(KEYINPUT57), .C1(new_n761_), .C2(new_n598_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n582_), .B1(new_n773_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n584_), .A2(new_n532_), .A3(new_n470_), .A4(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n781_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n470_), .A2(new_n565_), .A3(new_n569_), .A4(new_n582_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n671_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT120), .B1(new_n780_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n774_), .A2(new_n775_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n777_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n774_), .A2(KEYINPUT118), .A3(new_n775_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n764_), .A2(new_n772_), .A3(new_n765_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n583_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT120), .ZN(new_n794_));
  INV_X1    g593(.A(new_n786_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n362_), .A2(new_n291_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n616_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n787_), .A2(new_n324_), .A3(new_n796_), .A4(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G113gat), .B1(new_n800_), .B2(new_n671_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n773_), .A2(new_n788_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n583_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n623_), .B1(new_n804_), .B2(new_n795_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n798_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n802_), .A2(G113gat), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n801_), .B1(new_n808_), .B2(new_n671_), .ZN(G1340gat));
  NAND2_X1  g608(.A1(new_n802_), .A2(new_n807_), .ZN(new_n810_));
  OAI21_X1  g609(.A(G120gat), .B1(new_n810_), .B2(new_n470_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n242_), .B1(new_n470_), .B2(KEYINPUT60), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n800_), .B(new_n812_), .C1(KEYINPUT60), .C2(new_n242_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1341gat));
  INV_X1    g613(.A(G127gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n799_), .B2(new_n583_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n583_), .A2(new_n815_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n810_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT121), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n816_), .C1(new_n810_), .C2(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1342gat));
  AOI21_X1  g622(.A(G134gat), .B1(new_n800_), .B2(new_n599_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n570_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n810_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(G134gat), .ZN(G1343gat));
  NAND4_X1  g626(.A1(new_n787_), .A2(new_n616_), .A3(new_n796_), .A4(new_n623_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n797_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n671_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT122), .B(G141gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1344gat));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n471_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT123), .B(G148gat), .Z(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(G1345gat));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n582_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT61), .B(G155gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  AOI21_X1  g637(.A(G162gat), .B1(new_n829_), .B2(new_n599_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n828_), .A2(new_n825_), .A3(new_n797_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(G162gat), .B2(new_n840_), .ZN(G1347gat));
  NOR3_X1   g640(.A1(new_n616_), .A2(new_n291_), .A3(new_n362_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n805_), .A2(new_n842_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n843_), .A2(new_n532_), .A3(new_n217_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n671_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT124), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n845_), .A2(KEYINPUT124), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n805_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G169gat), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n849_), .A2(KEYINPUT62), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(KEYINPUT62), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n844_), .B1(new_n850_), .B2(new_n851_), .ZN(G1348gat));
  INV_X1    g651(.A(new_n843_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G176gat), .B1(new_n853_), .B2(new_n471_), .ZN(new_n854_));
  AND4_X1   g653(.A1(new_n324_), .A2(new_n787_), .A3(new_n796_), .A4(new_n842_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n471_), .A2(G176gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1349gat));
  AOI21_X1  g656(.A(G183gat), .B1(new_n855_), .B2(new_n582_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n843_), .A2(new_n212_), .A3(new_n583_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1350gat));
  OAI21_X1  g659(.A(G190gat), .B1(new_n843_), .B2(new_n825_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n599_), .A2(new_n213_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n843_), .B2(new_n862_), .ZN(G1351gat));
  NOR2_X1   g662(.A1(new_n362_), .A2(new_n291_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n828_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n671_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n471_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n871_), .A2(KEYINPUT126), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(KEYINPUT126), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n583_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT125), .Z(new_n876_));
  NAND2_X1  g675(.A1(new_n866_), .A2(new_n876_), .ZN(new_n877_));
  MUX2_X1   g676(.A(new_n872_), .B(new_n874_), .S(new_n877_), .Z(G1354gat));
  INV_X1    g677(.A(G218gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n866_), .B2(new_n570_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n599_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n828_), .A2(G218gat), .A3(new_n881_), .A4(new_n865_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n880_), .A2(KEYINPUT127), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT127), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n787_), .A2(new_n623_), .A3(new_n796_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n885_), .A2(new_n616_), .A3(new_n570_), .A4(new_n864_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G218gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n866_), .A2(new_n879_), .A3(new_n599_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n883_), .A2(new_n889_), .ZN(G1355gat));
endmodule


