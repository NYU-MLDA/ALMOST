//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n204_));
  OAI211_X1 g003(.A(new_n203_), .B(new_n204_), .C1(G155gat), .C2(G162gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n205_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(KEYINPUT3), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n206_), .A2(new_n211_), .A3(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G155gat), .B(G162gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT88), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n222_), .A3(new_n219_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n210_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT28), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G22gat), .B(G50gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n227_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n210_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n223_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n222_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT29), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT90), .B1(new_n224_), .B2(new_n225_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G197gat), .B(G204gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT21), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OR3_X1    g042(.A1(new_n238_), .A2(new_n242_), .A3(new_n239_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n237_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G228gat), .A2(G233gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT91), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n251_), .A3(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n234_), .A2(KEYINPUT29), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n253_), .A2(KEYINPUT89), .A3(new_n245_), .A4(new_n247_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(new_n252_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G78gat), .B(G106gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n230_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(KEYINPUT92), .Z(new_n262_));
  NAND4_X1  g061(.A1(new_n250_), .A2(new_n262_), .A3(new_n258_), .A4(new_n252_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT93), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n246_), .A2(new_n251_), .A3(new_n248_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n251_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n262_), .A4(new_n258_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n261_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n262_), .B1(new_n267_), .B2(new_n258_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n263_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n230_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275_));
  XOR2_X1   g074(.A(G8gat), .B(G36gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(G92gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT18), .B(G64gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT94), .ZN(new_n280_));
  OR2_X1    g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n285_));
  OAI211_X1 g084(.A(KEYINPUT24), .B(new_n281_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n281_), .A2(KEYINPUT24), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT23), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(new_n289_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT22), .B(G169gat), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n282_), .B(new_n283_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n291_), .B(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n296_), .B(new_n297_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT78), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n243_), .A2(new_n244_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT20), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n281_), .A2(KEYINPUT24), .A3(new_n282_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n289_), .A2(new_n292_), .A3(new_n290_), .A4(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n301_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n245_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n280_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  AOI211_X1 g116(.A(KEYINPUT94), .B(new_n317_), .C1(new_n307_), .C2(new_n312_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n303_), .A2(new_n305_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n308_), .B1(new_n320_), .B2(new_n245_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n245_), .A2(new_n311_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n279_), .B1(new_n319_), .B2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n293_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n304_), .B1(new_n293_), .B2(new_n301_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n245_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n245_), .A2(new_n311_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT20), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n315_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT94), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n313_), .A2(new_n280_), .A3(new_n315_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n323_), .A4(new_n279_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n275_), .B1(new_n324_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT98), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n279_), .B(KEYINPUT96), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n313_), .A2(new_n315_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n333_), .A2(new_n340_), .A3(KEYINPUT27), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT97), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n333_), .A2(new_n340_), .A3(KEYINPUT97), .A4(KEYINPUT27), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT84), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n234_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n224_), .A2(new_n351_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n348_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT4), .B1(new_n234_), .B2(new_n352_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n347_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n353_), .A2(new_n346_), .A3(new_n354_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT0), .B(G57gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT98), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n367_), .B(new_n275_), .C1(new_n324_), .C2(new_n334_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n336_), .A2(new_n345_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n352_), .B(KEYINPUT31), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n320_), .B(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G15gat), .B(G43gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT82), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n379_), .B(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n375_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n374_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n274_), .A2(new_n369_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n274_), .A2(new_n369_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n394_), .A3(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n363_), .A2(KEYINPUT33), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n357_), .A2(new_n358_), .A3(new_n398_), .A4(new_n362_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n346_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT95), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n362_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n353_), .A2(new_n347_), .A3(new_n354_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT95), .B(new_n346_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n324_), .A2(new_n334_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n400_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n319_), .A2(new_n323_), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n338_), .A2(new_n339_), .ZN(new_n412_));
  OAI221_X1 g211(.A(new_n411_), .B1(new_n412_), .B2(new_n410_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n270_), .A2(new_n273_), .A3(new_n409_), .A4(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n392_), .A2(new_n396_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT99), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT99), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n392_), .A2(new_n417_), .A3(new_n396_), .A4(new_n414_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n391_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G230gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G99gat), .A2(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT66), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(KEYINPUT6), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT66), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n422_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT67), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT7), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(G99gat), .C2(G106gat), .ZN(new_n430_));
  INV_X1    g229(.A(G99gat), .ZN(new_n431_));
  INV_X1    g230(.A(G106gat), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n431_), .B(new_n432_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n425_), .A2(KEYINPUT66), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n423_), .A2(KEYINPUT6), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(G99gat), .A4(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n427_), .A2(new_n434_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(G85gat), .A2(G92gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT68), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n444_), .A3(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT69), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n439_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(KEYINPUT8), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT10), .B(G99gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT64), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n431_), .A2(KEYINPUT10), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n431_), .A2(KEYINPUT10), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT64), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n432_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT65), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n441_), .A2(KEYINPUT9), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n432_), .C1(new_n454_), .C2(new_n457_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n440_), .A2(KEYINPUT9), .A3(new_n441_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n427_), .A2(new_n463_), .A3(new_n437_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n459_), .A2(new_n460_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n447_), .A2(KEYINPUT69), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n451_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT70), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n470_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT11), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n475_), .A3(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G71gat), .B(G78gat), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n473_), .B2(KEYINPUT11), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n468_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n480_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(new_n465_), .A3(new_n451_), .A4(new_n467_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(KEYINPUT12), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n468_), .A2(new_n487_), .A3(new_n482_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n421_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n420_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT71), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(KEYINPUT71), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT5), .B(G176gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G120gat), .B(G148gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n492_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT13), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(KEYINPUT72), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G29gat), .B(G36gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT15), .Z(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G1gat), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT75), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n516_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n524_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(KEYINPUT76), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n528_), .A2(new_n524_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n532_), .B1(new_n535_), .B2(new_n531_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n536_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n509_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT35), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n468_), .A2(new_n517_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(KEYINPUT73), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n552_), .B1(new_n516_), .B2(new_n468_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n553_), .B2(new_n549_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n547_), .B(new_n550_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT37), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n524_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n484_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n566_));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n571_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n565_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n573_), .B2(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n559_), .A2(KEYINPUT37), .A3(new_n560_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n562_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n419_), .A2(new_n542_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n366_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n519_), .A3(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT100), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT38), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n542_), .B(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n559_), .A2(new_n560_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(new_n576_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n416_), .A2(new_n418_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n391_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n587_), .A2(new_n590_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n366_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n583_), .A2(new_n584_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n585_), .A2(new_n596_), .A3(new_n597_), .ZN(G1324gat));
  AND2_X1   g397(.A1(new_n336_), .A2(new_n368_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(new_n345_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n580_), .A2(new_n520_), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n595_), .B2(new_n600_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n602_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n602_), .B(new_n607_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1325gat));
  OAI21_X1  g410(.A(G15gat), .B1(new_n595_), .B2(new_n396_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT103), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT103), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT41), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(KEYINPUT41), .A3(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n396_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n580_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n617_), .B(new_n618_), .C1(G15gat), .C2(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(G22gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n274_), .B(KEYINPUT104), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n594_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT42), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n622_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT105), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n580_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(G1327gat));
  NOR2_X1   g428(.A1(new_n419_), .A2(new_n542_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n588_), .A2(new_n577_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n366_), .A2(G29gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT107), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n578_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n561_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT43), .B1(new_n593_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n419_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n587_), .A4(new_n576_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n593_), .A2(KEYINPUT43), .A3(new_n638_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n419_), .B2(new_n637_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n587_), .A4(new_n576_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n581_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(G29gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n649_), .B2(G29gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n635_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  XNOR2_X1  g453(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(G36gat), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n630_), .A2(new_n657_), .A3(new_n601_), .A4(new_n631_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n600_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n643_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n662_), .B2(G36gat), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n656_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n657_), .B1(new_n661_), .B2(new_n643_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT108), .B(new_n655_), .C1(new_n666_), .C2(new_n660_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n643_), .A2(G43gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n648_), .A2(new_n389_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n632_), .A2(new_n619_), .ZN(new_n671_));
  OAI22_X1  g470(.A1(new_n669_), .A2(new_n670_), .B1(G43gat), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g472(.A(G50gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n623_), .A2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT110), .Z(new_n676_));
  NAND2_X1  g475(.A1(new_n632_), .A2(new_n676_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n643_), .A2(new_n274_), .A3(new_n648_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n674_), .ZN(G1331gat));
  NOR2_X1   g478(.A1(new_n419_), .A2(new_n541_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n579_), .A2(new_n509_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT111), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT111), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n581_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n509_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n680_), .A2(new_n687_), .A3(new_n590_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n581_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n686_), .B1(G57gat), .B2(new_n689_), .ZN(G1332gat));
  INV_X1    g489(.A(G64gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n685_), .A2(new_n691_), .A3(new_n601_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n688_), .B2(new_n601_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n694_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n685_), .A2(new_n698_), .A3(new_n619_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n688_), .B2(new_n619_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT49), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1334gat));
  INV_X1    g503(.A(G78gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n688_), .B2(new_n623_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n623_), .A2(new_n705_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT113), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n708_), .A2(new_n709_), .B1(new_n684_), .B2(new_n711_), .ZN(G1335gat));
  NOR2_X1   g511(.A1(new_n509_), .A2(new_n541_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n644_), .A2(new_n645_), .A3(new_n576_), .A4(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n581_), .A2(G85gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT115), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n680_), .A2(new_n687_), .A3(new_n631_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n720_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n366_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n718_), .B1(new_n723_), .B2(G85gat), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT116), .Z(G1336gat));
  AOI21_X1  g524(.A(new_n600_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n726_), .A2(KEYINPUT117), .A3(G92gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT117), .B1(new_n726_), .B2(G92gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n714_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n601_), .A2(G92gat), .ZN(new_n730_));
  AOI22_X1  g529(.A1(new_n727_), .A2(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(G1337gat));
  NAND2_X1  g530(.A1(new_n721_), .A2(new_n722_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n389_), .C1(new_n454_), .C2(new_n457_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G99gat), .B1(new_n714_), .B2(new_n396_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT51), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n732_), .A2(new_n432_), .A3(new_n274_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n729_), .A2(new_n274_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G106gat), .ZN(new_n743_));
  INV_X1    g542(.A(new_n274_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n741_), .B(G106gat), .C1(new_n714_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n740_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT53), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n740_), .B(new_n749_), .C1(new_n743_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1339gat));
  NOR2_X1   g550(.A1(new_n540_), .A2(new_n499_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n486_), .A2(new_n488_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n420_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n486_), .A2(new_n421_), .A3(new_n488_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n489_), .A2(KEYINPUT55), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n496_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n754_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n761_), .C2(new_n496_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT55), .B1(new_n755_), .B2(new_n420_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n757_), .B(new_n421_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n497_), .B1(new_n770_), .B2(new_n759_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n767_), .B1(new_n771_), .B2(KEYINPUT56), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n761_), .A2(new_n767_), .A3(KEYINPUT56), .A4(new_n496_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n753_), .B1(new_n766_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n531_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n530_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n539_), .B(new_n778_), .C1(new_n535_), .C2(new_n777_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT120), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n536_), .A2(new_n539_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(KEYINPUT120), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n501_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT57), .B(new_n588_), .C1(new_n776_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT118), .B1(new_n771_), .B2(KEYINPUT56), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n496_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT119), .ZN(new_n789_));
  INV_X1    g588(.A(new_n759_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n768_), .A2(new_n769_), .A3(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n754_), .B(new_n763_), .C1(new_n791_), .C2(new_n497_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n787_), .A2(new_n789_), .A3(new_n773_), .A4(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n784_), .B1(new_n793_), .B2(new_n752_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n786_), .B1(new_n794_), .B2(new_n589_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n762_), .A2(new_n763_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n788_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n783_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n498_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n797_), .A2(KEYINPUT58), .A3(new_n498_), .A4(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n638_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n785_), .A2(new_n795_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n576_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n636_), .A2(new_n561_), .A3(new_n576_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n541_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n601_), .A2(new_n366_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n389_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n744_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n274_), .B1(new_n805_), .B2(new_n812_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n816_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(KEYINPUT121), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n820_), .B1(new_n819_), .B2(new_n816_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n811_), .B1(new_n804_), .B2(new_n576_), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n825_), .A2(KEYINPUT59), .A3(new_n274_), .A4(new_n815_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT122), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n830_));
  OAI21_X1  g629(.A(G113gat), .B1(new_n540_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n822_), .A2(new_n827_), .A3(new_n829_), .A4(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n817_), .B2(new_n540_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1340gat));
  NAND3_X1  g633(.A1(new_n818_), .A2(new_n687_), .A3(new_n821_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT123), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n818_), .A2(new_n837_), .A3(new_n687_), .A4(new_n821_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(G120gat), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n817_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n509_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n840_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n843_), .ZN(G1341gat));
  NAND4_X1  g643(.A1(new_n822_), .A2(new_n827_), .A3(G127gat), .A4(new_n577_), .ZN(new_n845_));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n817_), .B2(new_n576_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n840_), .B2(new_n589_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n822_), .A2(new_n827_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT124), .B(G134gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n637_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n850_), .B2(new_n852_), .ZN(G1343gat));
  NAND3_X1  g652(.A1(new_n814_), .A2(new_n396_), .A3(new_n274_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT125), .Z(new_n855_));
  NOR2_X1   g654(.A1(new_n825_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n541_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n687_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n577_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n856_), .B2(new_n589_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n825_), .A2(new_n855_), .A3(new_n637_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(G162gat), .B2(new_n865_), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n600_), .A2(new_n581_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n619_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n623_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n813_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G169gat), .B1(new_n870_), .B2(new_n540_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n870_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n541_), .A3(new_n294_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT62), .B(G169gat), .C1(new_n870_), .C2(new_n540_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n873_), .A2(KEYINPUT126), .A3(new_n875_), .A4(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1348gat));
  AOI21_X1  g680(.A(G176gat), .B1(new_n874_), .B2(new_n687_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n825_), .A2(new_n274_), .A3(new_n868_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n509_), .A2(new_n295_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  NOR3_X1   g684(.A1(new_n870_), .A2(new_n576_), .A3(new_n287_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G183gat), .B1(new_n883_), .B2(new_n577_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n874_), .A2(new_n589_), .A3(new_n288_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G190gat), .B1(new_n870_), .B2(new_n637_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1351gat));
  NOR3_X1   g690(.A1(new_n825_), .A2(new_n619_), .A3(new_n744_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n867_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n540_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT127), .B(G197gat), .Z(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1352gat));
  INV_X1    g695(.A(new_n893_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n687_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g698(.A(KEYINPUT63), .B(G211gat), .C1(new_n897_), .C2(new_n577_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT63), .B(G211gat), .Z(new_n901_));
  AND3_X1   g700(.A1(new_n897_), .A2(new_n577_), .A3(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1354gat));
  NOR2_X1   g702(.A1(new_n893_), .A2(new_n588_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n897_), .A2(new_n638_), .ZN(new_n905_));
  MUX2_X1   g704(.A(new_n904_), .B(new_n905_), .S(G218gat), .Z(G1355gat));
endmodule


