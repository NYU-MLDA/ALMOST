//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n213_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT79), .B1(new_n213_), .B2(KEYINPUT23), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n212_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n210_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(KEYINPUT80), .A3(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G169gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n225_), .A3(new_n206_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT81), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n226_), .A2(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n225_), .A3(KEYINPUT81), .A4(new_n206_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(new_n212_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT82), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n221_), .A2(new_n222_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n212_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n213_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n220_), .B1(new_n242_), .B2(new_n217_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n210_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n222_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n233_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n233_), .A2(new_n246_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n247_), .A2(new_n229_), .A3(new_n228_), .A4(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  INV_X1    g050(.A(G99gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n237_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G15gat), .B(G43gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT83), .ZN(new_n256_));
  INV_X1    g055(.A(G71gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n259_));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n258_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n237_), .A2(new_n253_), .A3(new_n262_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT86), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT86), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n268_), .A3(new_n265_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT31), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n269_), .A2(new_n273_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G1gat), .B(G29gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT96), .B(G85gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G57gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G225gat), .A2(G233gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(G155gat), .B(G162gat), .Z(new_n284_));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n288_), .A2(new_n289_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(new_n287_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT87), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n297_), .B(new_n298_), .C1(new_n291_), .C2(KEYINPUT2), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n284_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n272_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(KEYINPUT4), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n300_), .A3(new_n272_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(KEYINPUT4), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT95), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT95), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n303_), .A2(new_n308_), .A3(KEYINPUT4), .A4(new_n305_), .ZN(new_n309_));
  AOI211_X1 g108(.A(new_n283_), .B(new_n304_), .C1(new_n307_), .C2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(new_n305_), .A3(new_n283_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n282_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n309_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n283_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n304_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n311_), .A3(new_n281_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n301_), .A2(KEYINPUT29), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT89), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  INV_X1    g125(.A(G218gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G211gat), .ZN(new_n328_));
  INV_X1    g127(.A(G211gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G218gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n326_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(G197gat), .A2(G204gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G197gat), .A2(G204gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT90), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  INV_X1    g134(.A(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n331_), .A2(new_n334_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n331_), .A2(new_n334_), .A3(new_n340_), .A4(KEYINPUT91), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n326_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(KEYINPUT21), .A3(new_n339_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT92), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n349_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n325_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n324_), .B1(new_n321_), .B2(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G78gat), .B(G106gat), .Z(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n363_));
  OR3_X1    g162(.A1(new_n301_), .A2(KEYINPUT29), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n301_), .B2(KEYINPUT29), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n359_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n356_), .A2(new_n370_), .A3(new_n357_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n360_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n360_), .B2(new_n371_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n352_), .A2(new_n355_), .A3(new_n250_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n208_), .B(KEYINPUT93), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n223_), .A2(new_n225_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n384_), .B2(new_n206_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n217_), .B1(new_n212_), .B2(new_n232_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n385_), .A2(new_n386_), .B1(new_n244_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n379_), .B1(new_n388_), .B2(new_n353_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n375_), .A2(new_n378_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n354_), .B1(new_n345_), .B2(new_n350_), .ZN(new_n391_));
  AOI211_X1 g190(.A(KEYINPUT92), .B(new_n349_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n235_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n385_), .A2(new_n386_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n244_), .A2(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n379_), .B1(new_n396_), .B2(new_n351_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n390_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT18), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n405_));
  INV_X1    g204(.A(new_n403_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n393_), .A2(new_n397_), .A3(new_n378_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n378_), .B1(new_n375_), .B2(new_n389_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AOI211_X1 g209(.A(KEYINPUT97), .B(new_n378_), .C1(new_n375_), .C2(new_n389_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n406_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT100), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT100), .B(new_n406_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n405_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n375_), .A2(new_n378_), .A3(new_n389_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT20), .B1(new_n388_), .B2(new_n353_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n352_), .A2(new_n355_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n235_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n417_), .B1(new_n420_), .B2(new_n378_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n406_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT27), .B1(new_n404_), .B2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n416_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n276_), .A2(new_n320_), .A3(new_n374_), .A4(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n318_), .B(new_n313_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n416_), .A2(new_n426_), .A3(new_n423_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n403_), .A2(KEYINPUT32), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT98), .B(new_n429_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n235_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT20), .B1(new_n396_), .B2(new_n351_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n377_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n433_), .A2(KEYINPUT97), .B1(new_n420_), .B2(new_n378_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n411_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n428_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n399_), .B2(new_n428_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n319_), .B(new_n430_), .C1(new_n436_), .C2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT99), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT98), .B1(new_n421_), .B2(new_n429_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT99), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n443_), .A2(new_n444_), .A3(new_n319_), .A4(new_n430_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n404_), .A2(new_n422_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n314_), .A2(new_n283_), .A3(new_n316_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n303_), .A2(new_n305_), .A3(new_n315_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n282_), .A3(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n318_), .A2(KEYINPUT33), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n318_), .A2(KEYINPUT33), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n446_), .B(new_n449_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n440_), .A2(new_n445_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n427_), .B1(new_n453_), .B2(new_n374_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n425_), .B1(new_n454_), .B2(new_n276_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G29gat), .B(G36gat), .Z(new_n456_));
  XOR2_X1   g255(.A(G43gat), .B(G50gat), .Z(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  INV_X1    g258(.A(G1gat), .ZN(new_n460_));
  INV_X1    g259(.A(G8gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G8gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n458_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n458_), .B(KEYINPUT15), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n465_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(new_n465_), .B2(new_n458_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(new_n468_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G113gat), .B(G141gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT78), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G169gat), .B(G197gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n473_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n455_), .A2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT67), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT6), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(new_n490_), .B2(new_n484_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n481_), .B(new_n482_), .C1(new_n487_), .C2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT8), .ZN(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT10), .B(G99gat), .Z(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT64), .B(G85gat), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n498_), .A2(G92gat), .B1(KEYINPUT9), .B2(new_n481_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT65), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n489_), .B(new_n496_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n493_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G78gat), .Z(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n503_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT12), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n493_), .A2(new_n510_), .A3(new_n502_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT69), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n517_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G120gat), .B(G148gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT5), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(KEYINPUT13), .A3(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n465_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n510_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G127gat), .B(G155gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n539_), .A2(KEYINPUT17), .A3(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n544_), .B(KEYINPUT17), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT76), .Z(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(KEYINPUT75), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n539_), .A2(KEYINPUT75), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n546_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT77), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n503_), .A2(new_n470_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT34), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n555_), .B(new_n560_), .C1(new_n458_), .C2(new_n503_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n559_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT71), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n555_), .B2(KEYINPUT72), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT36), .Z(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(KEYINPUT36), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(new_n573_), .A3(new_n566_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n572_), .A2(new_n576_), .A3(KEYINPUT37), .A4(new_n574_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n554_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n535_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n480_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n460_), .A3(new_n319_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT101), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n455_), .A2(new_n575_), .ZN(new_n588_));
  NOR4_X1   g387(.A1(new_n588_), .A2(new_n478_), .A3(new_n535_), .A4(new_n552_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n460_), .B1(new_n589_), .B2(new_n319_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n585_), .B2(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(G1324gat));
  INV_X1    g391(.A(new_n424_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n461_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT39), .Z(new_n595_));
  NAND3_X1  g394(.A1(new_n583_), .A2(new_n461_), .A3(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(G1325gat));
  INV_X1    g398(.A(G15gat), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n589_), .B2(new_n276_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT103), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT41), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT41), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n583_), .A2(new_n600_), .A3(new_n276_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(G1326gat));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n374_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n589_), .B2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT42), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n583_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1327gat));
  NAND3_X1  g411(.A1(new_n553_), .A2(new_n574_), .A3(new_n572_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT107), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(new_n535_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n480_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(G29gat), .B1(new_n617_), .B2(new_n319_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT43), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n579_), .A2(new_n580_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n453_), .A2(new_n374_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n427_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n276_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n274_), .A2(new_n275_), .ZN(new_n624_));
  NOR4_X1   g423(.A1(new_n593_), .A2(new_n624_), .A3(new_n319_), .A4(new_n608_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n619_), .B(new_n620_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n455_), .A2(KEYINPUT104), .A3(new_n619_), .A4(new_n620_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n455_), .A2(new_n620_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT43), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n535_), .A2(new_n478_), .A3(new_n554_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(KEYINPUT105), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT105), .B1(new_n632_), .B2(new_n633_), .ZN(new_n636_));
  NOR4_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(KEYINPUT106), .A4(KEYINPUT44), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n633_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT105), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n641_), .B2(new_n634_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT44), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(G29gat), .A3(new_n319_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n618_), .B1(new_n643_), .B2(new_n646_), .ZN(G1328gat));
  OAI211_X1 g446(.A(new_n593_), .B(new_n645_), .C1(new_n637_), .C2(new_n642_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G36gat), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT46), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT108), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n616_), .A2(G36gat), .A3(new_n424_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT45), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(KEYINPUT108), .B2(new_n650_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n649_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n649_), .B2(new_n654_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1329gat));
  XNOR2_X1  g456(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n276_), .A2(G43gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n644_), .B2(KEYINPUT44), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n637_), .B2(new_n642_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT109), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n660_), .B(new_n663_), .C1(new_n637_), .C2(new_n642_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G43gat), .B1(new_n617_), .B2(new_n276_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n658_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n658_), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n666_), .B(new_n669_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1330gat));
  AOI21_X1  g470(.A(G50gat), .B1(new_n617_), .B2(new_n608_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n645_), .A2(G50gat), .A3(new_n608_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n643_), .B2(new_n673_), .ZN(G1331gat));
  INV_X1    g473(.A(new_n535_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n581_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT111), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n455_), .A2(new_n478_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G57gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n319_), .ZN(new_n681_));
  NOR4_X1   g480(.A1(new_n588_), .A2(new_n675_), .A3(new_n479_), .A4(new_n553_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G57gat), .B1(new_n683_), .B2(new_n320_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1332gat));
  INV_X1    g484(.A(G64gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n682_), .B2(new_n593_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT48), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n679_), .A2(new_n686_), .A3(new_n593_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1333gat));
  AOI21_X1  g489(.A(new_n257_), .B1(new_n682_), .B2(new_n276_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT49), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n679_), .A2(new_n257_), .A3(new_n276_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1334gat));
  INV_X1    g493(.A(G78gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n682_), .B2(new_n608_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT50), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n679_), .A2(new_n695_), .A3(new_n608_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1335gat));
  NOR2_X1   g498(.A1(new_n614_), .A2(new_n675_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n678_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT112), .ZN(new_n702_));
  AOI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n319_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n675_), .A2(new_n479_), .A3(new_n554_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n632_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n320_), .A2(new_n497_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(G1336gat));
  AOI21_X1  g506(.A(G92gat), .B1(new_n702_), .B2(new_n593_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n593_), .A2(G92gat), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT113), .Z(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n705_), .B2(new_n710_), .ZN(G1337gat));
  AND2_X1   g510(.A1(new_n276_), .A2(new_n494_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT114), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n702_), .A2(new_n712_), .B1(new_n713_), .B2(KEYINPUT51), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n705_), .A2(new_n276_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n252_), .B2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n713_), .A2(KEYINPUT51), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n716_), .B(new_n717_), .Z(G1338gat));
  NAND3_X1  g517(.A1(new_n702_), .A2(new_n495_), .A3(new_n608_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT116), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n705_), .A2(new_n608_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G106gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n720_), .A3(G106gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g527(.A(G113gat), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT117), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n529_), .A2(new_n730_), .A3(new_n479_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n520_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT117), .B1(new_n732_), .B2(new_n478_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n520_), .A2(KEYINPUT55), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n517_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n516_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n515_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n520_), .B2(KEYINPUT55), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n527_), .B1(new_n736_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT56), .B(new_n527_), .C1(new_n736_), .C2(new_n740_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n734_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n477_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n473_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n467_), .B1(new_n472_), .B2(KEYINPUT118), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(KEYINPUT118), .B2(new_n472_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n477_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n531_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n531_), .A2(KEYINPUT119), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n575_), .B1(new_n745_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n529_), .A2(new_n751_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n761_), .A2(KEYINPUT58), .B1(new_n579_), .B2(new_n580_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n743_), .A2(new_n744_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n760_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT57), .B(new_n575_), .C1(new_n745_), .C2(new_n756_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n759_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n552_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n582_), .A2(new_n478_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(KEYINPUT54), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(KEYINPUT54), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n276_), .A2(new_n319_), .A3(new_n374_), .A4(new_n424_), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT120), .Z(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n729_), .B1(new_n776_), .B2(new_n478_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT121), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n771_), .A2(new_n772_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n768_), .B2(new_n553_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n775_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(KEYINPUT59), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT122), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n779_), .B1(new_n768_), .B2(new_n552_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT59), .B1(new_n785_), .B2(new_n781_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT122), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n757_), .A2(new_n758_), .B1(new_n762_), .B2(new_n765_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n554_), .B1(new_n788_), .B2(new_n767_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n787_), .B(new_n782_), .C1(new_n789_), .C2(new_n779_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n784_), .A2(new_n786_), .A3(new_n790_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n791_), .A2(new_n729_), .A3(new_n478_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n777_), .A2(KEYINPUT121), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n778_), .A2(new_n792_), .A3(new_n793_), .ZN(G1340gat));
  NAND4_X1  g593(.A1(new_n784_), .A2(new_n786_), .A3(new_n535_), .A4(new_n790_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G120gat), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT60), .ZN(new_n797_));
  AOI21_X1  g596(.A(G120gat), .B1(new_n535_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n797_), .B2(G120gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n773_), .A2(new_n775_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n796_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT123), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n796_), .A2(KEYINPUT123), .A3(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1341gat));
  OAI21_X1  g604(.A(G127gat), .B1(new_n791_), .B2(new_n552_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n553_), .A2(G127gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n776_), .B2(new_n807_), .ZN(G1342gat));
  OR3_X1    g607(.A1(new_n776_), .A2(G134gat), .A3(new_n575_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n791_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n810_));
  INV_X1    g609(.A(G134gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(G1343gat));
  NOR4_X1   g611(.A1(new_n276_), .A2(new_n593_), .A3(new_n320_), .A4(new_n374_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n773_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n478_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(new_n288_), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n675_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n289_), .ZN(G1345gat));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n814_), .B2(new_n553_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n773_), .A2(KEYINPUT124), .A3(new_n554_), .A4(new_n813_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1346gat));
  AOI21_X1  g623(.A(new_n814_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n825_));
  INV_X1    g624(.A(G162gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n572_), .A2(new_n826_), .A3(new_n574_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n825_), .A2(new_n826_), .B1(new_n814_), .B2(new_n827_), .ZN(G1347gat));
  NOR3_X1   g627(.A1(new_n624_), .A2(new_n424_), .A3(new_n319_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n780_), .A2(new_n608_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n205_), .B1(new_n831_), .B2(new_n479_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(KEYINPUT62), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n479_), .A3(new_n384_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(KEYINPUT62), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(G1348gat));
  AOI21_X1  g635(.A(G176gat), .B1(new_n831_), .B2(new_n535_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n785_), .A2(new_n608_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n675_), .A2(new_n206_), .A3(new_n830_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(G1349gat));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n554_), .A3(new_n829_), .ZN(new_n841_));
  INV_X1    g640(.A(G183gat), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n552_), .A2(new_n202_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n841_), .A2(new_n842_), .B1(new_n831_), .B2(new_n843_), .ZN(G1350gat));
  NAND4_X1  g643(.A1(new_n831_), .A2(new_n203_), .A3(new_n574_), .A4(new_n572_), .ZN(new_n845_));
  INV_X1    g644(.A(G190gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n831_), .B2(new_n620_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n848_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n849_), .B2(new_n850_), .ZN(G1351gat));
  NOR3_X1   g650(.A1(new_n276_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n773_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n479_), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n854_), .A2(KEYINPUT126), .A3(new_n335_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT126), .B1(new_n854_), .B2(new_n335_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n335_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(G1352gat));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n535_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n859_), .B(new_n860_), .Z(G1353gat));
  INV_X1    g660(.A(new_n552_), .ZN(new_n862_));
  AOI211_X1 g661(.A(KEYINPUT63), .B(G211gat), .C1(new_n853_), .C2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n853_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n552_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT63), .B(G211gat), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n865_), .B2(new_n866_), .ZN(G1354gat));
  AND2_X1   g666(.A1(new_n853_), .A2(new_n620_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n572_), .A2(new_n327_), .A3(new_n574_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n868_), .A2(new_n327_), .B1(new_n864_), .B2(new_n869_), .ZN(G1355gat));
endmodule


