//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G197gat), .B(G204gat), .Z(new_n208_));
  OR2_X1    g007(.A1(new_n208_), .A2(KEYINPUT21), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(KEYINPUT21), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n217_), .A2(KEYINPUT24), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT78), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(G183gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT78), .B1(new_n231_), .B2(KEYINPUT25), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n222_), .B(new_n227_), .C1(new_n229_), .C2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT82), .B1(new_n223_), .B2(KEYINPUT23), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT22), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT22), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n220_), .A2(KEYINPUT80), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G176gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n241_), .A2(new_n243_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT81), .A3(new_n217_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n239_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT81), .B1(new_n247_), .B2(new_n217_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n234_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT83), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n234_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n215_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n228_), .A2(new_n230_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n222_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n237_), .A2(new_n238_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT80), .B(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT22), .B(G169gat), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n260_), .A2(new_n261_), .B1(G169gat), .B2(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT89), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n227_), .A2(new_n235_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n262_), .B2(KEYINPUT89), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n259_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT20), .B1(new_n267_), .B2(new_n214_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G226gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT19), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n255_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n252_), .A2(new_n254_), .A3(new_n215_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n267_), .B2(new_n214_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n207_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n254_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n247_), .A2(new_n217_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT81), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n248_), .A3(new_n239_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n253_), .B1(new_n282_), .B2(new_n234_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n214_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n266_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n285_), .A2(new_n263_), .B1(new_n258_), .B2(new_n257_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n274_), .B1(new_n286_), .B2(new_n215_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n287_), .A3(new_n272_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n273_), .A2(new_n275_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n206_), .B(new_n288_), .C1(new_n289_), .C2(new_n272_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT27), .B1(new_n277_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n273_), .A2(new_n272_), .A3(new_n275_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n272_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n207_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT98), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n270_), .B1(new_n255_), .B2(new_n268_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n292_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT98), .A3(new_n207_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT27), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n271_), .A2(new_n276_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n206_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n291_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G57gat), .B(G85gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT94), .ZN(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G29gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  NOR2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT84), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G155gat), .A3(G162gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n312_), .B1(new_n317_), .B2(KEYINPUT1), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n314_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT85), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n314_), .A2(new_n316_), .A3(new_n322_), .A4(new_n319_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G141gat), .B(G148gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327_));
  INV_X1    g126(.A(G141gat), .ZN(new_n328_));
  INV_X1    g127(.A(G148gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n330_), .A2(new_n333_), .A3(new_n334_), .A4(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n312_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n326_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G127gat), .B(G134gat), .Z(new_n341_));
  XOR2_X1   g140(.A(G113gat), .B(G120gat), .Z(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT90), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT86), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n326_), .B2(new_n339_), .ZN(new_n346_));
  AOI211_X1 g145(.A(KEYINPUT86), .B(new_n338_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n344_), .B1(new_n348_), .B2(new_n343_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  NOR4_X1   g149(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT90), .A4(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT4), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n340_), .A2(KEYINPUT86), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n338_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n345_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT92), .B(KEYINPUT4), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n353_), .A2(new_n355_), .A3(new_n343_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT91), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n352_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n353_), .A2(new_n364_), .A3(new_n355_), .A4(new_n343_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(new_n344_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n359_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n311_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n361_), .B1(new_n367_), .B2(KEYINPUT4), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n353_), .A2(new_n355_), .A3(new_n343_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n364_), .B1(new_n354_), .B2(new_n350_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n373_), .A2(new_n365_), .B1(G225gat), .B2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n311_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n370_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT97), .B1(new_n369_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT97), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n373_), .B2(new_n365_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n368_), .B(new_n311_), .C1(new_n381_), .C2(new_n361_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n305_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT28), .B1(new_n348_), .B2(KEYINPUT29), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n386_), .B(new_n387_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G22gat), .B(G50gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n385_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G228gat), .ZN(new_n395_));
  INV_X1    g194(.A(G233gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n214_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n348_), .B2(KEYINPUT29), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n214_), .B1(new_n354_), .B2(new_n387_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n395_), .A2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT88), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n346_), .A2(new_n347_), .A3(new_n387_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n405_), .B(new_n401_), .C1(new_n406_), .C2(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT87), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n404_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n394_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n403_), .A2(new_n407_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n404_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n414_), .A2(KEYINPUT87), .A3(new_n408_), .A4(new_n393_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G43gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n252_), .A2(new_n418_), .A3(new_n254_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n420_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT31), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n420_), .A2(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT31), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n420_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n428_), .A2(new_n434_), .A3(new_n343_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n343_), .B1(new_n428_), .B2(new_n434_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n416_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n426_), .A2(new_n427_), .A3(KEYINPUT31), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n432_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n350_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n428_), .A2(new_n434_), .A3(new_n343_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n411_), .A2(new_n443_), .A3(new_n415_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n384_), .B1(new_n438_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n298_), .B2(new_n292_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n303_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n369_), .B2(new_n376_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT95), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n376_), .A2(new_n451_), .A3(KEYINPUT33), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n277_), .A2(new_n290_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n382_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n358_), .A2(new_n359_), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n381_), .A2(KEYINPUT96), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT96), .B1(new_n381_), .B2(new_n456_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n311_), .B1(new_n367_), .B2(new_n360_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT95), .B1(new_n382_), .B2(new_n454_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n452_), .A2(new_n455_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n446_), .B1(new_n450_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n445_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G232gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT34), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G29gat), .B(G36gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n467_), .A2(KEYINPUT68), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(KEYINPUT68), .ZN(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  OR3_X1    g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT15), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G85gat), .B(G92gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT9), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(KEYINPUT10), .B(G99gat), .Z(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n479_), .A2(new_n480_), .A3(G85gat), .A4(G92gat), .ZN(new_n487_));
  AND3_X1   g286(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n483_), .A2(new_n486_), .A3(new_n487_), .A4(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n485_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT65), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n497_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n492_), .B1(new_n505_), .B2(new_n478_), .ZN(new_n506_));
  AOI211_X1 g305(.A(KEYINPUT8), .B(new_n477_), .C1(new_n497_), .C2(new_n490_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n491_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n475_), .A2(new_n476_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n476_), .B1(new_n475_), .B2(new_n508_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n497_), .A2(new_n490_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n492_), .A3(new_n478_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT65), .B1(new_n500_), .B2(new_n501_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n495_), .A2(new_n496_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n477_), .B1(new_n516_), .B2(new_n502_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n517_), .B2(new_n492_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT66), .B1(new_n518_), .B2(new_n491_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT66), .B(new_n491_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n519_), .A2(new_n521_), .A3(new_n473_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT35), .B(new_n466_), .C1(new_n511_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n510_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n475_), .A2(new_n476_), .A3(new_n508_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n466_), .A2(KEYINPUT35), .ZN(new_n527_));
  INV_X1    g326(.A(new_n522_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n466_), .A2(KEYINPUT35), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT36), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n523_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n533_), .B(KEYINPUT36), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n464_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G78gat), .Z(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n543_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n508_), .A2(KEYINPUT12), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT66), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n508_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n551_), .B2(new_n520_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n552_), .B2(KEYINPUT12), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n520_), .A3(new_n547_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT67), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n553_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n548_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n555_), .B1(new_n561_), .B2(new_n554_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NOR3_X1   g365(.A1(new_n560_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(KEYINPUT13), .A3(new_n569_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n473_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G15gat), .B(G22gat), .ZN(new_n576_));
  INV_X1    g375(.A(G8gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G8gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  NAND3_X1  g380(.A1(new_n575_), .A2(KEYINPUT75), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n581_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n473_), .A2(new_n474_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT15), .B1(new_n471_), .B2(new_n472_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT76), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT76), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n586_), .A2(new_n590_), .A3(new_n595_), .A4(new_n592_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n582_), .A2(new_n585_), .B1(new_n473_), .B2(new_n587_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n594_), .B(new_n596_), .C1(new_n592_), .C2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT77), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(KEYINPUT77), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n574_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n547_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT70), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(new_n581_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n581_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n619_), .A2(KEYINPUT71), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT71), .B1(new_n619_), .B2(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n615_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n620_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT74), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n619_), .A2(KEYINPUT74), .A3(new_n620_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n613_), .B(KEYINPUT17), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n608_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n540_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n377_), .A2(new_n383_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n202_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT99), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT37), .B1(new_n535_), .B2(new_n538_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT37), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n523_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n523_), .A2(new_n530_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n637_), .B(new_n638_), .C1(new_n639_), .C2(new_n537_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n630_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n464_), .A2(new_n608_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n202_), .A3(new_n633_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT38), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n635_), .A2(new_n646_), .ZN(G1324gat));
  AOI21_X1  g446(.A(KEYINPUT98), .B1(new_n299_), .B2(new_n207_), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n296_), .B(new_n206_), .C1(new_n298_), .C2(new_n292_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n304_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n291_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n577_), .B1(new_n632_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n644_), .A2(new_n577_), .A3(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  AOI21_X1  g458(.A(new_n422_), .B1(new_n632_), .B2(new_n443_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT100), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n644_), .A2(new_n422_), .A3(new_n443_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT101), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n540_), .A2(new_n631_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n416_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G22gat), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n644_), .A2(new_n672_), .A3(new_n416_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT102), .Z(G1327gat));
  NAND4_X1  g474(.A1(new_n607_), .A2(new_n572_), .A3(new_n630_), .A4(new_n573_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n539_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n379_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n652_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n411_), .A2(new_n443_), .A3(new_n415_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n443_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n462_), .A2(new_n450_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n446_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n678_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n678_), .A2(new_n688_), .A3(KEYINPUT104), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n633_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n636_), .A2(new_n640_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n695_), .B(new_n696_), .C1(new_n445_), .C2(new_n463_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT103), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n445_), .B2(new_n463_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT43), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n688_), .A2(new_n701_), .A3(new_n695_), .A4(new_n696_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n676_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n703_), .B2(new_n704_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n633_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n694_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NOR2_X1   g508(.A1(new_n305_), .A2(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n691_), .A2(new_n692_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n714_));
  NAND4_X1  g513(.A1(new_n691_), .A2(KEYINPUT106), .A3(new_n692_), .A4(new_n710_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n713_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n703_), .A2(new_n704_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G36gat), .B1(new_n723_), .B2(new_n305_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n718_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n718_), .B2(new_n724_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NAND2_X1  g527(.A1(new_n693_), .A2(new_n443_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT109), .B(G43gat), .Z(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n443_), .A2(G43gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT108), .B1(new_n707_), .B2(new_n733_), .ZN(new_n734_));
  AND4_X1   g533(.A1(KEYINPUT108), .A2(new_n721_), .A3(new_n722_), .A4(new_n733_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n731_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n693_), .B2(new_n416_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n416_), .A2(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n707_), .B2(new_n742_), .ZN(G1331gat));
  NOR4_X1   g542(.A1(new_n464_), .A2(new_n643_), .A3(new_n607_), .A4(new_n574_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n633_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n574_), .A2(new_n630_), .A3(new_n607_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n540_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n633_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(KEYINPUT110), .ZN(new_n750_));
  MUX2_X1   g549(.A(KEYINPUT110), .B(new_n750_), .S(G57gat), .Z(new_n751_));
  AOI21_X1  g550(.A(new_n745_), .B1(new_n748_), .B2(new_n751_), .ZN(G1332gat));
  OAI21_X1  g551(.A(G64gat), .B1(new_n747_), .B2(new_n305_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n744_), .A2(new_n756_), .A3(new_n652_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n747_), .B2(new_n437_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  INV_X1    g560(.A(G71gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n744_), .A2(new_n762_), .A3(new_n443_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n747_), .B2(new_n669_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  INV_X1    g565(.A(G78gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n744_), .A2(new_n767_), .A3(new_n416_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n464_), .A2(new_n607_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n572_), .A2(new_n573_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n630_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n677_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n633_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT113), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n772_), .A2(new_n607_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n703_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(G85gat), .A3(new_n633_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1336gat));
  INV_X1    g580(.A(G92gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n775_), .A2(new_n782_), .A3(new_n652_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n779_), .A2(new_n652_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n782_), .ZN(G1337gat));
  NAND2_X1  g584(.A1(new_n443_), .A2(new_n484_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n779_), .A2(new_n443_), .ZN(new_n787_));
  OAI221_X1 g586(.A(KEYINPUT114), .B1(new_n774_), .B2(new_n786_), .C1(new_n787_), .C2(new_n494_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n775_), .A2(new_n485_), .A3(new_n416_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n779_), .A2(new_n416_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G106gat), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT52), .B(new_n485_), .C1(new_n779_), .C2(new_n416_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n790_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n603_), .B1(new_n597_), .B2(new_n593_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n586_), .A2(new_n593_), .A3(new_n590_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n804_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n554_), .B(new_n549_), .C1(new_n552_), .C2(KEYINPUT12), .ZN(new_n811_));
  INV_X1    g610(.A(new_n555_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n560_), .B2(KEYINPUT55), .ZN(new_n814_));
  INV_X1    g613(.A(new_n549_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT12), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n561_), .B2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n554_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n558_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n817_), .B(KEYINPUT55), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT56), .B(new_n566_), .C1(new_n814_), .C2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT117), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n820_), .A3(new_n813_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT117), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n566_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n566_), .B1(new_n814_), .B2(new_n821_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n829_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n823_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n604_), .A2(new_n605_), .A3(new_n568_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n810_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n802_), .B1(new_n837_), .B2(new_n539_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n809_), .A2(new_n567_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n822_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n566_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n641_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n839_), .B(KEYINPUT58), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n566_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n830_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n824_), .A2(new_n825_), .B1(new_n812_), .B2(new_n811_), .ZN(new_n849_));
  AOI211_X1 g648(.A(new_n847_), .B(new_n848_), .C1(new_n849_), .C2(new_n820_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n829_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n827_), .B2(new_n566_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n835_), .B1(new_n853_), .B2(new_n823_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n677_), .C1(new_n854_), .C2(new_n810_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n838_), .A2(new_n846_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n630_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n574_), .A2(new_n606_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n643_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n771_), .A2(new_n607_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n858_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n861_), .A2(new_n642_), .A3(new_n641_), .A4(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n749_), .B1(new_n857_), .B2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n444_), .A2(new_n652_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n801_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n856_), .B2(new_n630_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n867_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n869_), .A2(new_n749_), .A3(new_n870_), .A4(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n800_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n866_), .A2(new_n867_), .A3(new_n871_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n869_), .A2(new_n749_), .A3(new_n870_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n875_), .B(KEYINPUT120), .C1(new_n801_), .C2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(G113gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n606_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(new_n877_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n876_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n881_), .B2(new_n606_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1340gat));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n574_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n876_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n884_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n868_), .A2(new_n873_), .A3(new_n574_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n884_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n630_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n874_), .A2(new_n877_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n881_), .B2(new_n630_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1342gat));
  INV_X1    g692(.A(G134gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n641_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n874_), .A2(new_n877_), .A3(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n881_), .B2(new_n677_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1343gat));
  NOR4_X1   g697(.A1(new_n869_), .A2(new_n749_), .A3(new_n438_), .A4(new_n652_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n607_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n771_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n642_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  INV_X1    g705(.A(G162gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n899_), .A2(new_n907_), .A3(new_n539_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n899_), .A2(new_n696_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n416_), .B1(new_n857_), .B2(new_n865_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n652_), .A2(new_n443_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n633_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n606_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n911_), .B1(new_n916_), .B2(new_n219_), .ZN(new_n917_));
  OAI211_X1 g716(.A(KEYINPUT62), .B(G169gat), .C1(new_n915_), .C2(new_n606_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n261_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(G1348gat));
  OAI21_X1  g719(.A(new_n677_), .B1(new_n854_), .B2(new_n810_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n921_), .A2(new_n802_), .B1(new_n845_), .B2(new_n844_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n642_), .B1(new_n922_), .B2(new_n855_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT121), .B(new_n669_), .C1(new_n923_), .C2(new_n864_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n869_), .B2(new_n416_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n914_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n928_), .A2(new_n574_), .A3(new_n220_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n912_), .A2(new_n771_), .A3(new_n914_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n927_), .A2(new_n929_), .B1(new_n260_), .B2(new_n930_), .ZN(G1349gat));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n630_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n924_), .A2(new_n926_), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n231_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n228_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(KEYINPUT122), .B1(new_n912_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939_));
  NOR4_X1   g738(.A1(new_n869_), .A2(new_n939_), .A3(new_n416_), .A4(new_n936_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n934_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n934_), .A2(new_n941_), .A3(KEYINPUT123), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n915_), .B2(new_n641_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n539_), .A2(new_n230_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n915_), .B2(new_n948_), .ZN(G1351gat));
  INV_X1    g748(.A(new_n869_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n438_), .A2(new_n633_), .A3(new_n305_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(G197gat), .ZN(new_n953_));
  OR4_X1    g752(.A1(KEYINPUT124), .A2(new_n952_), .A3(new_n953_), .A4(new_n606_), .ZN(new_n954_));
  AND2_X1   g753(.A1(new_n950_), .A2(new_n951_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n607_), .ZN(new_n956_));
  OAI21_X1  g755(.A(KEYINPUT124), .B1(new_n956_), .B2(new_n953_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n953_), .ZN(new_n958_));
  AND3_X1   g757(.A1(new_n954_), .A2(new_n957_), .A3(new_n958_), .ZN(G1352gat));
  NOR2_X1   g758(.A1(new_n952_), .A2(new_n574_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(KEYINPUT125), .B(G204gat), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1353gat));
  NOR2_X1   g761(.A1(new_n952_), .A2(new_n630_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964_));
  XOR2_X1   g763(.A(KEYINPUT63), .B(G211gat), .Z(new_n965_));
  AND3_X1   g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n963_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n964_), .B1(new_n963_), .B2(new_n965_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n966_), .A2(new_n967_), .A3(new_n968_), .ZN(G1354gat));
  INV_X1    g768(.A(G218gat), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n955_), .A2(new_n970_), .A3(new_n539_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n952_), .A2(new_n641_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(new_n970_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(KEYINPUT127), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n971_), .B(new_n975_), .C1(new_n970_), .C2(new_n972_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1355gat));
endmodule


