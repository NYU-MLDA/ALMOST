//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204_));
  OR4_X1    g003(.A1(new_n204_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n205_));
  OAI22_X1  g004(.A1(new_n204_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT8), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n211_), .A3(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT10), .B(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n219_), .B(new_n223_), .C1(new_n208_), .C2(new_n220_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n218_), .A2(new_n224_), .A3(new_n203_), .A4(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n213_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n228_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G232gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT35), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT15), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n234_), .B(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT72), .B1(new_n227_), .B2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n235_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n239_), .A2(new_n240_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G134gat), .B(G162gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  INV_X1    g049(.A(KEYINPUT36), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n245_), .A2(new_n246_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n247_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n250_), .B(KEYINPUT36), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n247_), .B2(new_n254_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT37), .B1(new_n255_), .B2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n245_), .B(new_n246_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n256_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT37), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n247_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G71gat), .B(G78gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G57gat), .B(G64gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT11), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT11), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n269_), .A2(new_n266_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G231gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275_));
  INV_X1    g074(.A(G1gat), .ZN(new_n276_));
  INV_X1    g075(.A(G8gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT14), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT73), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n274_), .B(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G155gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G183gat), .B(G211gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n289_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n283_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n291_), .B2(new_n283_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n265_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G230gat), .A2(G233gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT64), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n272_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n227_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n272_), .B1(new_n213_), .B2(new_n226_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n299_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT68), .ZN(new_n304_));
  NOR2_X1   g103(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n213_), .A2(new_n226_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n306_), .B2(new_n272_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n227_), .A2(new_n300_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n302_), .A2(KEYINPUT69), .A3(KEYINPUT12), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n307_), .A2(new_n310_), .A3(new_n298_), .A4(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(new_n299_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n304_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G176gat), .B(G204gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(G120gat), .B(G148gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n304_), .A2(new_n312_), .A3(new_n314_), .A4(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(KEYINPUT13), .A3(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n296_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(KEYINPUT75), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(KEYINPUT75), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n281_), .A2(new_n234_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n243_), .B2(new_n281_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G229gat), .A2(G233gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n281_), .A2(new_n234_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G113gat), .B(G141gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT76), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G169gat), .B(G197gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(new_n338_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352_));
  INV_X1    g151(.A(G141gat), .ZN(new_n353_));
  INV_X1    g152(.A(G148gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT85), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT2), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(KEYINPUT85), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n357_), .A2(new_n360_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n355_), .A2(new_n356_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n351_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n369_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n350_), .A2(KEYINPUT1), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G155gat), .A3(G162gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n376_), .A3(new_n349_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n353_), .A2(new_n354_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n358_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n366_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n371_), .A2(new_n381_), .A3(new_n372_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n367_), .A2(new_n369_), .A3(KEYINPUT82), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n379_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n363_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n356_), .B2(new_n355_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n355_), .A2(new_n356_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n360_), .A4(new_n362_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n389_), .B2(new_n351_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n380_), .B(KEYINPUT4), .C1(new_n384_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n366_), .A2(new_n379_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n382_), .A2(new_n383_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n391_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n395_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n401_), .A2(new_n380_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n392_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n391_), .A2(KEYINPUT89), .A3(new_n393_), .A4(new_n397_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  NAND4_X1  g207(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n409_), .A2(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(KEYINPUT33), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n393_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n408_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n391_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT26), .B(G190gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT25), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G183gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT77), .B(G183gat), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n417_), .B(new_n419_), .C1(new_n420_), .C2(new_n418_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422_));
  INV_X1    g221(.A(G169gat), .ZN(new_n423_));
  INV_X1    g222(.A(G176gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT78), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n423_), .A2(new_n424_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G169gat), .A2(G176gat), .ZN(new_n433_));
  OR3_X1    g232(.A1(new_n432_), .A2(new_n422_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n425_), .A2(new_n428_), .A3(new_n435_), .A4(new_n429_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n421_), .A2(new_n431_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT22), .B(G169gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n438_), .B2(new_n424_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n420_), .A2(G190gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n428_), .A2(new_n429_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT79), .ZN(new_n444_));
  XOR2_X1   g243(.A(G197gat), .B(G204gat), .Z(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT21), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G197gat), .B(G204gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT21), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G211gat), .B(G218gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  OR3_X1    g250(.A1(new_n447_), .A2(new_n450_), .A3(new_n448_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n437_), .A2(new_n454_), .A3(new_n442_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n444_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n430_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT25), .B(G183gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n417_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n434_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n439_), .B1(new_n441_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n451_), .A2(new_n452_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(KEYINPUT20), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G226gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT19), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(new_n222_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT18), .B(G64gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n437_), .A2(new_n454_), .A3(new_n442_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n454_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n464_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n468_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT20), .B1(new_n463_), .B2(new_n464_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n469_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n473_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT88), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n469_), .A2(new_n480_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n473_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n469_), .A2(new_n480_), .A3(new_n473_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n412_), .A2(new_n416_), .A3(new_n483_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT90), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n473_), .A2(KEYINPUT32), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n484_), .B2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n469_), .A2(KEYINPUT90), .A3(new_n492_), .A4(new_n480_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n476_), .A2(new_n479_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(new_n468_), .ZN(new_n499_));
  AOI211_X1 g298(.A(KEYINPUT91), .B(new_n477_), .C1(new_n476_), .C2(new_n479_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n456_), .A2(KEYINPUT20), .A3(new_n477_), .A4(new_n465_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n492_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n468_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT91), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n497_), .A3(new_n468_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT92), .B1(new_n509_), .B2(new_n493_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n496_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n414_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n409_), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n512_), .A2(new_n514_), .A3(new_n414_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n490_), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n519_));
  NAND2_X1  g318(.A1(G227gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G71gat), .B(G99gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(KEYINPUT81), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n524_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n444_), .A2(KEYINPUT81), .A3(new_n455_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G43gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n528_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n523_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n474_), .A2(new_n475_), .A3(new_n524_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT81), .B1(new_n444_), .B2(new_n455_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n527_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n523_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n529_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n384_), .B(KEYINPUT31), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT83), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n532_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT83), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT87), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G78gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n546_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n453_), .B1(new_n394_), .B2(KEYINPUT29), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n217_), .B1(new_n390_), .B2(new_n552_), .ZN(new_n553_));
  AND4_X1   g352(.A1(new_n552_), .A2(new_n366_), .A3(new_n217_), .A4(new_n379_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n551_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(G106gat), .B1(new_n394_), .B2(KEYINPUT29), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n464_), .B1(new_n390_), .B2(new_n552_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n390_), .A2(new_n552_), .A3(new_n217_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G22gat), .B(G50gat), .Z(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n555_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n550_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n555_), .A2(new_n559_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n560_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n555_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n549_), .A3(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n544_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n568_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n532_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n530_), .A2(new_n531_), .A3(new_n523_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n536_), .B1(new_n535_), .B2(new_n529_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n572_), .B(new_n573_), .C1(new_n576_), .C2(new_n542_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n571_), .A2(new_n577_), .B1(new_n516_), .B2(new_n515_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT27), .B1(new_n486_), .B2(new_n488_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n473_), .B(KEYINPUT94), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n481_), .B1(new_n509_), .B2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n581_), .B2(KEYINPUT27), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n518_), .A2(new_n570_), .B1(new_n578_), .B2(new_n582_), .ZN(new_n583_));
  NOR4_X1   g382(.A1(new_n330_), .A2(new_n331_), .A3(new_n348_), .A4(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n517_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT38), .B1(new_n586_), .B2(new_n276_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n261_), .A2(new_n263_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n583_), .A2(new_n591_), .A3(new_n294_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n328_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n592_), .A2(new_n347_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n276_), .B1(new_n594_), .B2(new_n585_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n586_), .A2(KEYINPUT38), .A3(new_n276_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT95), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n586_), .A2(new_n598_), .A3(KEYINPUT38), .A4(new_n276_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n589_), .A2(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(new_n582_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n584_), .A2(new_n277_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n594_), .A2(new_n602_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n605_), .B2(G8gat), .ZN(new_n606_));
  AOI211_X1 g405(.A(KEYINPUT39), .B(new_n277_), .C1(new_n594_), .C2(new_n602_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g408(.A(G15gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n594_), .B2(new_n544_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT41), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n584_), .A2(new_n610_), .A3(new_n544_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1326gat));
  INV_X1    g413(.A(G22gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n594_), .B2(new_n569_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT42), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n584_), .A2(new_n615_), .A3(new_n569_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1327gat));
  NAND4_X1  g418(.A1(new_n326_), .A2(new_n347_), .A3(new_n327_), .A4(new_n294_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n583_), .A2(KEYINPUT43), .A3(new_n265_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n571_), .A2(new_n577_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n517_), .A3(new_n582_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n504_), .B1(new_n503_), .B2(new_n492_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n509_), .A2(KEYINPUT92), .A3(new_n493_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n626_), .A2(new_n627_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n483_), .A2(new_n489_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n416_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n628_), .A2(new_n585_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n570_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n625_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n265_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n623_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n621_), .B1(new_n622_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n621_), .B(new_n641_), .C1(new_n622_), .C2(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n517_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n583_), .A2(new_n590_), .A3(new_n620_), .ZN(new_n645_));
  INV_X1    g444(.A(G29gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n585_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(G1328gat));
  INV_X1    g447(.A(KEYINPUT46), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n640_), .A2(new_n602_), .A3(new_n642_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G36gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G36gat), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT45), .ZN(new_n655_));
  INV_X1    g454(.A(G36gat), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n582_), .B(KEYINPUT99), .Z(new_n657_));
  NAND4_X1  g456(.A1(new_n645_), .A2(KEYINPUT101), .A3(new_n656_), .A4(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n634_), .A2(new_n656_), .A3(new_n621_), .A4(new_n591_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n657_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n658_), .A2(new_n659_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n659_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n655_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT100), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n659_), .A3(new_n663_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(KEYINPUT45), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n649_), .B1(new_n654_), .B2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n666_), .A2(new_n670_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(KEYINPUT46), .C1(new_n653_), .C2(new_n652_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1329gat));
  AND2_X1   g474(.A1(new_n645_), .A2(new_n544_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(G43gat), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n640_), .A2(G43gat), .A3(new_n544_), .A4(new_n642_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n678_), .A2(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT47), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n677_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n643_), .B2(new_n572_), .ZN(new_n687_));
  INV_X1    g486(.A(G50gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n645_), .A2(new_n688_), .A3(new_n569_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1331gat));
  INV_X1    g489(.A(G57gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n294_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n348_), .A3(new_n328_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n583_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT103), .Z(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n695_), .B2(new_n517_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n592_), .A2(new_n348_), .A3(new_n328_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(new_n691_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n517_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT104), .Z(G1332gat));
  OAI21_X1  g499(.A(G64gat), .B1(new_n697_), .B2(new_n662_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT48), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n662_), .A2(G64gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n695_), .B2(new_n703_), .ZN(G1333gat));
  INV_X1    g503(.A(new_n544_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n697_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G71gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G71gat), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n695_), .A2(new_n705_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n711_), .B(new_n712_), .C1(G71gat), .C2(new_n713_), .ZN(G1334gat));
  OAI21_X1  g513(.A(G78gat), .B1(new_n697_), .B2(new_n572_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT50), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n572_), .A2(G78gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n695_), .B2(new_n717_), .ZN(G1335gat));
  NAND3_X1  g517(.A1(new_n328_), .A2(new_n348_), .A3(new_n294_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n583_), .A2(new_n719_), .A3(new_n590_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G85gat), .B1(new_n720_), .B2(new_n585_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT43), .B1(new_n583_), .B2(new_n265_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n634_), .A2(new_n623_), .A3(new_n635_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(new_n221_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n721_), .B1(new_n726_), .B2(new_n585_), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n720_), .B2(new_n602_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n725_), .A2(new_n222_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n657_), .ZN(G1337gat));
  NAND3_X1  g529(.A1(new_n720_), .A2(new_n216_), .A3(new_n544_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT106), .ZN(new_n732_));
  OAI21_X1  g531(.A(G99gat), .B1(new_n725_), .B2(new_n705_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT108), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n734_), .A2(KEYINPUT107), .A3(KEYINPUT108), .A4(KEYINPUT51), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n734_), .A2(KEYINPUT107), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(G1338gat));
  AOI21_X1  g539(.A(new_n217_), .B1(new_n724_), .B2(new_n569_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n744_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n720_), .A2(new_n217_), .A3(new_n569_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT53), .B1(new_n748_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n747_), .A2(new_n753_), .A3(new_n749_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  INV_X1    g554(.A(G113gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n323_), .A2(new_n347_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n323_), .A2(KEYINPUT111), .A3(new_n347_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n307_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n299_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n312_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n763_), .A2(new_n762_), .A3(new_n299_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n320_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n302_), .B(new_n309_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n298_), .B1(new_n771_), .B2(new_n307_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n312_), .B1(new_n772_), .B2(new_n762_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n767_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n320_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n761_), .B1(new_n770_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n333_), .A2(new_n336_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n334_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n343_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n346_), .A2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT112), .Z(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n324_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n590_), .B1(new_n777_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n782_), .A2(new_n323_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n320_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n769_), .B(new_n322_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n787_), .B(KEYINPUT58), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n635_), .A3(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT57), .B(new_n590_), .C1(new_n777_), .C2(new_n783_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n786_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n294_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n692_), .A2(new_n348_), .A3(new_n327_), .A4(new_n326_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n797_), .A2(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n602_), .A2(new_n517_), .A3(new_n577_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n756_), .B1(new_n804_), .B2(new_n348_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT113), .B(new_n756_), .C1(new_n804_), .C2(new_n348_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(new_n795_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n786_), .A2(new_n794_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(KEYINPUT115), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n786_), .A2(new_n794_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n295_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n803_), .B(new_n810_), .C1(new_n816_), .C2(new_n800_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n804_), .A2(KEYINPUT59), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT116), .B(G113gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n348_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n809_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  XNOR2_X1  g621(.A(KEYINPUT117), .B(G120gat), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT60), .B1(new_n328_), .B2(new_n824_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n804_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(KEYINPUT60), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n826_), .A2(new_n817_), .A3(new_n328_), .A4(new_n818_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n804_), .B2(new_n294_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT118), .B(new_n830_), .C1(new_n804_), .C2(new_n294_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n294_), .A2(new_n830_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n819_), .B2(new_n836_), .ZN(G1342gat));
  NAND4_X1  g636(.A1(new_n817_), .A2(new_n818_), .A3(G134gat), .A4(new_n635_), .ZN(new_n838_));
  INV_X1    g637(.A(G134gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n804_), .B2(new_n590_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1343gat));
  AOI21_X1  g640(.A(new_n800_), .B1(new_n796_), .B2(new_n294_), .ZN(new_n842_));
  NOR4_X1   g641(.A1(new_n842_), .A2(new_n517_), .A3(new_n571_), .A4(new_n657_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n347_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n328_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n850_), .A3(new_n295_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n843_), .B2(new_n295_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n853_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1346gat));
  NOR2_X1   g656(.A1(new_n842_), .A2(new_n571_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n585_), .A3(new_n662_), .ZN(new_n859_));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n265_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n859_), .B2(new_n590_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT120), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(new_n860_), .C1(new_n859_), .C2(new_n590_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n863_), .B2(new_n865_), .ZN(G1347gat));
  XNOR2_X1  g665(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(KEYINPUT122), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n657_), .A2(new_n517_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n577_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n816_), .B2(new_n800_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n348_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n423_), .B1(new_n867_), .B2(KEYINPUT122), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n868_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n438_), .ZN(new_n876_));
  OAI221_X1 g675(.A(new_n873_), .B1(KEYINPUT122), .B2(new_n867_), .C1(new_n871_), .C2(new_n348_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  NAND2_X1  g677(.A1(new_n802_), .A2(new_n870_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n879_), .A2(new_n424_), .A3(new_n593_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n871_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n328_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n882_), .B2(new_n424_), .ZN(G1349gat));
  INV_X1    g682(.A(new_n458_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n881_), .A2(KEYINPUT123), .A3(new_n884_), .A4(new_n295_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n420_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n879_), .B2(new_n294_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n295_), .B(new_n870_), .C1(new_n816_), .C2(new_n800_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n458_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n885_), .A2(new_n887_), .A3(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n871_), .B2(new_n265_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n591_), .A2(new_n417_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT124), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n871_), .B2(new_n894_), .ZN(G1351gat));
  NOR4_X1   g694(.A1(new_n842_), .A2(new_n348_), .A3(new_n571_), .A4(new_n869_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT126), .B1(new_n896_), .B2(KEYINPUT125), .ZN(new_n897_));
  AOI21_X1  g696(.A(G197gat), .B1(new_n896_), .B2(KEYINPUT125), .ZN(new_n898_));
  INV_X1    g697(.A(new_n571_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n869_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n802_), .A2(new_n347_), .A3(new_n899_), .A4(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n897_), .A2(new_n898_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n898_), .B1(new_n897_), .B2(new_n904_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1352gat));
  NAND2_X1  g706(.A1(new_n858_), .A2(new_n900_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n593_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(new_n910_), .ZN(G1353gat));
  NOR2_X1   g712(.A1(new_n908_), .A2(new_n294_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AND2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  INV_X1    g717(.A(G218gat), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n908_), .A2(new_n919_), .A3(new_n265_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n858_), .A2(new_n591_), .A3(new_n900_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(new_n921_), .ZN(G1355gat));
endmodule


