//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n576_,
    new_n577_, new_n578_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT15), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT76), .ZN(new_n209_));
  INV_X1    g008(.A(G15gat), .ZN(new_n210_));
  INV_X1    g009(.A(G22gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G15gat), .A2(G22gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G1gat), .A2(G8gat), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n212_), .A2(new_n213_), .B1(KEYINPUT14), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n209_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n206_), .A2(KEYINPUT15), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n207_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n206_), .A2(new_n216_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT78), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n206_), .A2(new_n216_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n219_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(KEYINPUT77), .A3(new_n223_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT78), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n218_), .A2(new_n230_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n222_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G141gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n222_), .A2(new_n229_), .A3(new_n231_), .A4(new_n235_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT23), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(KEYINPUT24), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT88), .ZN(new_n246_));
  INV_X1    g045(.A(G169gat), .ZN(new_n247_));
  INV_X1    g046(.A(G176gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT24), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n249_), .A2(new_n250_), .A3(new_n243_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n242_), .B1(G183gat), .B2(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n249_), .B1(new_n256_), .B2(new_n248_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n246_), .A2(new_n254_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G197gat), .B(G204gat), .Z(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(KEYINPUT21), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(KEYINPUT21), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n261_), .A2(new_n262_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT20), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n256_), .A2(KEYINPUT81), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n247_), .A2(KEYINPUT22), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n248_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OAI221_X1 g071(.A(new_n255_), .B1(new_n247_), .B2(new_n248_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n274_));
  NOR2_X1   g073(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n275_));
  OAI21_X1  g074(.A(G190gat), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT80), .ZN(new_n277_));
  INV_X1    g076(.A(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT26), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(new_n252_), .A3(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n245_), .A2(new_n251_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n273_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n268_), .B1(new_n265_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT19), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n282_), .A2(new_n265_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n287_), .B(KEYINPUT20), .C1(new_n266_), .C2(new_n258_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n285_), .B(KEYINPUT87), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G8gat), .B(G36gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n286_), .A2(new_n298_), .A3(new_n290_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(KEYINPUT90), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT90), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n291_), .A2(new_n302_), .A3(new_n296_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n283_), .A2(new_n285_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n288_), .A2(new_n289_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(KEYINPUT27), .B(new_n299_), .C1(new_n307_), .C2(new_n298_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT3), .Z(new_n316_));
  NAND2_X1  g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT2), .Z(new_n318_));
  OAI211_X1 g117(.A(new_n313_), .B(new_n314_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n314_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n313_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n315_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n317_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n265_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G233gat), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n328_), .A2(KEYINPUT85), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(KEYINPUT85), .ZN(new_n330_));
  OAI21_X1  g129(.A(G228gat), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G78gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G106gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G22gat), .B(G50gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n336_), .B(G106gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n325_), .A2(new_n326_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT28), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n331_), .A2(new_n332_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G15gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n282_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G134gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G113gat), .B(G120gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n355_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  INV_X1    g159(.A(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n359_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n325_), .B(new_n358_), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT4), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n325_), .A2(KEYINPUT4), .A3(new_n358_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  INV_X1    g172(.A(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n368_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n369_), .A2(new_n378_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n372_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(KEYINPUT94), .A3(new_n381_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n367_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n310_), .A2(new_n352_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT95), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT95), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n310_), .A2(new_n352_), .A3(new_n389_), .A4(new_n386_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n350_), .A2(new_n351_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n300_), .A2(new_n303_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT91), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n370_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n377_), .B1(new_n369_), .B2(new_n378_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n395_), .A2(KEYINPUT93), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT93), .B1(new_n395_), .B2(new_n396_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  OAI22_X1  g198(.A1(new_n397_), .A2(new_n398_), .B1(new_n381_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n381_), .A2(new_n399_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n381_), .A2(KEYINPUT92), .A3(new_n399_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n400_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n300_), .A2(new_n406_), .A3(new_n303_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n394_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n298_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n286_), .A2(new_n409_), .A3(new_n290_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n382_), .B(new_n410_), .C1(new_n409_), .C2(new_n307_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n392_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n384_), .A2(new_n385_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n352_), .A2(new_n309_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n367_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n240_), .B1(new_n391_), .B2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT10), .B(G99gat), .Z(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n337_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G85gat), .B(G92gat), .Z(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT9), .ZN(new_n420_));
  INV_X1    g219(.A(G92gat), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n374_), .A2(new_n421_), .A3(KEYINPUT9), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G99gat), .A2(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT6), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(G99gat), .A3(G106gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n418_), .A2(new_n420_), .A3(new_n422_), .A4(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n429_));
  NOR2_X1   g228(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n430_));
  OAI22_X1  g229(.A1(new_n429_), .A2(new_n430_), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n432_));
  INV_X1    g231(.A(G99gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n337_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n427_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT8), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n419_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n425_), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n423_), .A2(KEYINPUT6), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT65), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n424_), .A2(new_n426_), .A3(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n441_), .A2(new_n443_), .A3(new_n431_), .A4(new_n434_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n437_), .B1(new_n444_), .B2(new_n419_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n438_), .B1(new_n445_), .B2(KEYINPUT66), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447_));
  AOI211_X1 g246(.A(new_n447_), .B(new_n437_), .C1(new_n444_), .C2(new_n419_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n428_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n217_), .A3(new_n207_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G232gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT34), .ZN(new_n452_));
  INV_X1    g251(.A(new_n428_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n419_), .ZN(new_n454_));
  AOI211_X1 g253(.A(KEYINPUT8), .B(new_n454_), .C1(new_n435_), .C2(new_n427_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n431_), .A2(new_n434_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n424_), .A2(new_n426_), .A3(new_n442_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n442_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT8), .B1(new_n459_), .B2(new_n454_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n455_), .B1(new_n460_), .B2(new_n447_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n448_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n453_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n206_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT74), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n449_), .A2(new_n466_), .A3(new_n206_), .ZN(new_n467_));
  OAI221_X1 g266(.A(new_n450_), .B1(KEYINPUT35), .B2(new_n452_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n452_), .A2(KEYINPUT35), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT71), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n468_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G190gat), .B(G218gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G134gat), .B(G162gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(KEYINPUT36), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(KEYINPUT36), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n471_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n479_), .B(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G57gat), .B(G64gat), .Z(new_n483_));
  INV_X1    g282(.A(KEYINPUT11), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT67), .B(G71gat), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n335_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT67), .B(G71gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G78gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT68), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n485_), .A2(new_n487_), .A3(new_n492_), .A4(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n483_), .A2(new_n484_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n216_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G127gat), .B(G155gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT16), .ZN(new_n504_));
  XOR2_X1   g303(.A(G183gat), .B(G211gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT17), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n502_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n482_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n497_), .A2(new_n498_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n463_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT12), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n449_), .A2(new_n517_), .A3(new_n499_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n449_), .B2(new_n499_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT69), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n463_), .A2(new_n515_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n449_), .A2(new_n499_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n514_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n516_), .B(new_n525_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n521_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT5), .ZN(new_n529_));
  XOR2_X1   g328(.A(G176gat), .B(G204gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(KEYINPUT70), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(KEYINPUT13), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n512_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n416_), .A2(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT96), .ZN(new_n542_));
  INV_X1    g341(.A(G1gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(KEYINPUT96), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n413_), .A4(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT38), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n479_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n391_), .B2(new_n415_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n539_), .A2(new_n240_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n511_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n413_), .ZN(new_n555_));
  OAI21_X1  g354(.A(G1gat), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(new_n546_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n556_), .A3(new_n557_), .ZN(G1324gat));
  INV_X1    g357(.A(G8gat), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n542_), .A2(new_n559_), .A3(new_n309_), .A4(new_n544_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT97), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n553_), .B2(new_n309_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT39), .Z(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n561_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(G1325gat));
  INV_X1    g366(.A(new_n367_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n210_), .B1(new_n553_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT99), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT41), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(KEYINPUT41), .ZN(new_n572_));
  INV_X1    g371(.A(new_n541_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n210_), .A3(new_n568_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(G1326gat));
  AOI21_X1  g374(.A(new_n211_), .B1(new_n553_), .B2(new_n392_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT42), .Z(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n211_), .A3(new_n392_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1327gat));
  INV_X1    g378(.A(G29gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n391_), .A2(new_n415_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n482_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(KEYINPUT100), .A3(KEYINPUT43), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT43), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n482_), .B1(new_n391_), .B2(new_n415_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n584_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n511_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n550_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT44), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT44), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n594_), .B(new_n591_), .C1(new_n584_), .C2(new_n588_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n580_), .B1(new_n596_), .B2(new_n413_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n539_), .A2(new_n511_), .A3(new_n479_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n416_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n413_), .A2(new_n580_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT101), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n597_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n598_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1328gat));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT46), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n611_));
  INV_X1    g410(.A(G36gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n596_), .B2(new_n309_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n600_), .A2(new_n612_), .A3(new_n309_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT45), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n610_), .B(new_n611_), .C1(new_n613_), .C2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n589_), .A2(new_n592_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n594_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n589_), .A2(KEYINPUT44), .A3(new_n592_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n309_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G36gat), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n622_), .A2(new_n608_), .A3(new_n609_), .A4(new_n615_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n617_), .A2(new_n623_), .ZN(G1329gat));
  AOI21_X1  g423(.A(G43gat), .B1(new_n600_), .B2(new_n568_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT104), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n619_), .A2(new_n620_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n568_), .A2(G43gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g429(.A(G50gat), .B1(new_n600_), .B2(new_n392_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n392_), .A2(G50gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n596_), .B2(new_n632_), .ZN(G1331gat));
  INV_X1    g432(.A(new_n539_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(new_n239_), .A3(new_n590_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n549_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G57gat), .B1(new_n637_), .B2(new_n555_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n634_), .A2(new_n239_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n581_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n512_), .ZN(new_n641_));
  INV_X1    g440(.A(G57gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n413_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(G1332gat));
  INV_X1    g443(.A(G64gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n636_), .B2(new_n309_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT48), .Z(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n645_), .A3(new_n309_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1333gat));
  INV_X1    g448(.A(G71gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n636_), .B2(new_n568_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT49), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n650_), .A3(new_n568_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1334gat));
  NAND3_X1  g453(.A1(new_n641_), .A2(new_n335_), .A3(new_n392_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G78gat), .B1(new_n637_), .B2(new_n352_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT106), .ZN(G1335gat));
  NAND2_X1  g461(.A1(new_n639_), .A2(new_n590_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G85gat), .B1(new_n665_), .B2(new_n555_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n640_), .A2(new_n511_), .A3(new_n479_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n374_), .A3(new_n413_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1336gat));
  OAI21_X1  g468(.A(G92gat), .B1(new_n665_), .B2(new_n310_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n667_), .A2(new_n421_), .A3(new_n309_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT107), .ZN(G1337gat));
  OAI21_X1  g472(.A(G99gat), .B1(new_n665_), .B2(new_n367_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n568_), .A3(new_n417_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g476(.A1(new_n667_), .A2(new_n337_), .A3(new_n392_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT52), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n664_), .A2(new_n392_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(G106gat), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT52), .B(new_n337_), .C1(new_n664_), .C2(new_n392_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g483(.A(KEYINPUT119), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n482_), .A2(new_n240_), .A3(new_n634_), .A4(new_n511_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT55), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n521_), .A2(new_n689_), .A3(new_n526_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n521_), .A2(KEYINPUT110), .A3(new_n689_), .A4(new_n526_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT12), .B1(new_n463_), .B2(new_n515_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n449_), .A2(new_n517_), .A3(new_n499_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n523_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT111), .B1(new_n697_), .B2(new_n513_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n518_), .A2(new_n519_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n699_), .B(new_n514_), .C1(new_n700_), .C2(new_n523_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n520_), .B2(new_n689_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n695_), .A2(new_n696_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n704_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n516_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n698_), .A2(new_n701_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n694_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT56), .A3(new_n534_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT115), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT116), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n533_), .B1(new_n694_), .B2(new_n706_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(KEYINPUT56), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT115), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n713_), .A3(KEYINPUT56), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT56), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n698_), .A2(new_n701_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n703_), .A2(new_n705_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT116), .B(new_n715_), .C1(new_n719_), .C2(new_n533_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n709_), .A2(new_n712_), .A3(new_n714_), .A4(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n226_), .A2(new_n219_), .A3(new_n228_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n218_), .A2(new_n227_), .A3(new_n220_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n236_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n238_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT113), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n532_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n721_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n721_), .B(new_n727_), .C1(KEYINPUT117), .C2(KEYINPUT58), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n582_), .A3(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n733_));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n532_), .A2(new_n734_), .A3(new_n239_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n532_), .B2(new_n239_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT56), .B1(new_n707_), .B2(new_n534_), .ZN(new_n738_));
  AOI211_X1 g537(.A(new_n715_), .B(new_n533_), .C1(new_n694_), .C2(new_n706_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n726_), .A2(new_n536_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n733_), .B1(new_n742_), .B2(new_n479_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n732_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT118), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n482_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n743_), .B1(new_n747_), .B2(new_n731_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT118), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n751_), .B(new_n548_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n746_), .A2(new_n750_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n688_), .B1(new_n754_), .B2(new_n590_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n310_), .A2(new_n352_), .A3(new_n413_), .A4(new_n568_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n756_), .A2(KEYINPUT59), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n685_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n752_), .B1(new_n745_), .B2(KEYINPUT118), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n511_), .B1(new_n760_), .B2(new_n750_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT119), .B(new_n757_), .C1(new_n761_), .C2(new_n688_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n748_), .A2(new_n753_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n688_), .B1(new_n763_), .B2(new_n590_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT59), .B1(new_n764_), .B2(new_n756_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n759_), .A2(new_n762_), .A3(new_n239_), .A4(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G113gat), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n764_), .A2(new_n756_), .ZN(new_n768_));
  INV_X1    g567(.A(G113gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n239_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1340gat));
  NAND4_X1  g570(.A1(new_n759_), .A2(new_n762_), .A3(new_n539_), .A4(new_n765_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G120gat), .ZN(new_n773_));
  INV_X1    g572(.A(G120gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n634_), .B2(KEYINPUT60), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n768_), .B(new_n775_), .C1(KEYINPUT60), .C2(new_n774_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1341gat));
  NAND4_X1  g576(.A1(new_n759_), .A2(new_n762_), .A3(new_n511_), .A4(new_n765_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G127gat), .ZN(new_n779_));
  INV_X1    g578(.A(G127gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n768_), .A2(new_n780_), .A3(new_n511_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1342gat));
  NAND4_X1  g581(.A1(new_n759_), .A2(new_n762_), .A3(new_n582_), .A4(new_n765_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G134gat), .ZN(new_n784_));
  INV_X1    g583(.A(G134gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n768_), .A2(new_n785_), .A3(new_n548_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1343gat));
  XOR2_X1   g586(.A(new_n686_), .B(new_n687_), .Z(new_n788_));
  AOI211_X1 g587(.A(new_n752_), .B(new_n743_), .C1(new_n747_), .C2(new_n731_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n511_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n555_), .A2(new_n352_), .A3(new_n309_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n367_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n239_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT120), .B(G141gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1344gat));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n539_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g596(.A(KEYINPUT61), .B(G155gat), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n792_), .A2(new_n800_), .A3(new_n511_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n792_), .B2(new_n511_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n803_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n801_), .A3(new_n798_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1346gat));
  NAND3_X1  g606(.A1(new_n792_), .A2(G162gat), .A3(new_n582_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n790_), .A2(new_n367_), .A3(new_n548_), .A4(new_n791_), .ZN(new_n809_));
  INV_X1    g608(.A(G162gat), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(KEYINPUT122), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT122), .B1(new_n809_), .B2(new_n810_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT123), .B(new_n808_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1347gat));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n352_), .A2(new_n309_), .A3(new_n386_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n753_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT118), .B(new_n743_), .C1(new_n747_), .C2(new_n731_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n590_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n240_), .B(new_n819_), .C1(new_n822_), .C2(new_n788_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n818_), .B1(new_n823_), .B2(new_n247_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n819_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n239_), .B(new_n825_), .C1(new_n761_), .C2(new_n688_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(KEYINPUT62), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n256_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT124), .B1(new_n826_), .B2(G169gat), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n828_), .A2(new_n833_), .ZN(G1348gat));
  NOR2_X1   g633(.A1(new_n755_), .A2(new_n819_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G176gat), .B1(new_n835_), .B2(new_n539_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n764_), .A2(new_n819_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n634_), .A2(new_n248_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1349gat));
  AOI21_X1  g638(.A(G183gat), .B1(new_n837_), .B2(new_n511_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n590_), .A2(new_n252_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n835_), .B2(new_n841_), .ZN(G1350gat));
  NAND2_X1  g641(.A1(new_n548_), .A2(new_n253_), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(KEYINPUT125), .Z(new_n844_));
  NAND2_X1  g643(.A1(new_n835_), .A2(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n755_), .A2(new_n482_), .A3(new_n819_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n278_), .ZN(G1351gat));
  NOR2_X1   g646(.A1(new_n764_), .A2(new_n568_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n310_), .A2(new_n352_), .A3(new_n413_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n240_), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n851_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n634_), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(G204gat), .Z(G1353gat));
  XOR2_X1   g653(.A(KEYINPUT63), .B(G211gat), .Z(new_n855_));
  NAND4_X1  g654(.A1(new_n848_), .A2(new_n511_), .A3(new_n849_), .A4(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT126), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n850_), .B2(new_n590_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n856_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n861_), .B2(KEYINPUT126), .ZN(G1354gat));
  INV_X1    g661(.A(G218gat), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n850_), .A2(new_n863_), .A3(new_n482_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n850_), .A2(KEYINPUT127), .A3(new_n479_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(G218gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT127), .B1(new_n850_), .B2(new_n479_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(G1355gat));
endmodule


