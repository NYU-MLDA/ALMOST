//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT78), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n210_), .B(new_n211_), .C1(G183gat), .C2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n203_), .A2(new_n214_), .A3(new_n204_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n206_), .A2(new_n212_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n217_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n204_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(new_n209_), .B2(KEYINPUT77), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G183gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n222_), .B(new_n225_), .C1(KEYINPUT76), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(KEYINPUT76), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n218_), .B(new_n221_), .C1(new_n228_), .C2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n216_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n216_), .A2(new_n232_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G43gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n243_), .B(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n202_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n241_), .A2(new_n202_), .A3(new_n246_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n235_), .A2(KEYINPUT80), .A3(new_n238_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT82), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT82), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n254_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(new_n255_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n250_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n250_), .A2(new_n264_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n248_), .A2(new_n249_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n249_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(new_n247_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT2), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(KEYINPUT84), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT85), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(KEYINPUT85), .B(new_n272_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT3), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .A4(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n286_), .B2(KEYINPUT1), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(KEYINPUT83), .A3(G155gat), .A4(G162gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n286_), .A2(KEYINPUT1), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .A4(new_n285_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n282_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n272_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n289_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT94), .B1(new_n258_), .B2(new_n259_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n297_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n284_), .B2(new_n288_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n262_), .A2(new_n255_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT94), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n257_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n299_), .A2(new_n306_), .A3(KEYINPUT4), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n298_), .A2(new_n260_), .A3(new_n310_), .A4(new_n263_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n307_), .B(KEYINPUT95), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n308_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G29gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G57gat), .B(G85gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n308_), .B(new_n319_), .C1(new_n309_), .C2(new_n313_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  XOR2_X1   g127(.A(G197gat), .B(G204gat), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT21), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G197gat), .B(G204gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT21), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G218gat), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n337_), .A2(G211gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(G211gat), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT86), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n330_), .B(new_n333_), .C1(new_n336_), .C2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT86), .B1(new_n338_), .B2(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n335_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT21), .A4(new_n329_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n328_), .B1(new_n236_), .B2(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n213_), .A2(KEYINPUT92), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n213_), .A2(KEYINPUT92), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n212_), .A2(new_n205_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  AND4_X1   g148(.A1(new_n210_), .A2(new_n221_), .A3(new_n211_), .A4(new_n217_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT26), .B(G190gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n230_), .A2(new_n227_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n230_), .B2(new_n227_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n355_), .A3(KEYINPUT91), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT91), .B1(new_n350_), .B2(new_n355_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n349_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n327_), .B(new_n346_), .C1(new_n359_), .C2(new_n345_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G8gat), .B(G36gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT18), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT20), .B1(new_n236_), .B2(new_n345_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n359_), .B2(new_n345_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n360_), .B(new_n364_), .C1(new_n366_), .C2(new_n327_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n341_), .A2(new_n344_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n328_), .B1(new_n233_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n349_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n358_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n356_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n371_), .B1(new_n374_), .B2(new_n370_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n326_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n376_), .A2(KEYINPUT97), .A3(new_n364_), .A4(new_n360_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT27), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n350_), .A2(new_n355_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n380_), .A3(new_n349_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n346_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n326_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n375_), .B2(new_n326_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n364_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n323_), .B1(new_n378_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n345_), .B1(new_n302_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G228gat), .ZN(new_n391_));
  INV_X1    g190(.A(G233gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  OAI221_X1 g193(.A(new_n345_), .B1(new_n391_), .B2(new_n392_), .C1(new_n302_), .C2(new_n389_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n289_), .A2(new_n389_), .A3(new_n297_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT28), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n302_), .A2(new_n400_), .A3(new_n389_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G22gat), .B(G50gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n397_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n396_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n388_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n399_), .A2(new_n401_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n402_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n403_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n409_), .A2(new_n413_), .A3(KEYINPUT87), .A4(new_n397_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n396_), .A2(KEYINPUT88), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n394_), .A2(new_n395_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n403_), .A3(new_n412_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n367_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n376_), .A2(KEYINPUT93), .A3(new_n364_), .A4(new_n360_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n360_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n359_), .A2(new_n345_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n327_), .B1(new_n427_), .B2(new_n371_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n385_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n425_), .A3(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n430_), .A2(KEYINPUT98), .A3(new_n379_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT98), .B1(new_n430_), .B2(new_n379_), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n387_), .B(new_n422_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n322_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n299_), .A2(new_n306_), .A3(KEYINPUT4), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT33), .A3(new_n308_), .A4(new_n319_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n299_), .A2(new_n306_), .A3(new_n312_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n320_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n435_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n322_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n319_), .B1(new_n437_), .B2(new_n308_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n384_), .A2(KEYINPUT32), .A3(new_n364_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n376_), .A2(new_n447_), .A3(new_n360_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n442_), .A2(new_n430_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n420_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n271_), .B1(new_n433_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n378_), .A2(new_n386_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n271_), .A2(new_n451_), .A3(new_n445_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G1gat), .ZN(new_n459_));
  INV_X1    g258(.A(G8gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT71), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT71), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(KEYINPUT14), .C1(new_n459_), .C2(new_n460_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G1gat), .B(G8gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n468_), .B(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n476_));
  INV_X1    g275(.A(new_n468_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n468_), .A2(new_n471_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n475_), .A2(new_n480_), .A3(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n458_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n492_));
  INV_X1    g291(.A(G231gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(new_n392_), .ZN(new_n494_));
  INV_X1    g293(.A(G64gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G57gat), .ZN(new_n496_));
  INV_X1    g295(.A(G57gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G64gat), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n496_), .A2(new_n498_), .A3(KEYINPUT64), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT64), .B1(new_n496_), .B2(new_n498_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT11), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(G64gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n495_), .A2(G57gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT11), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n496_), .A2(new_n498_), .A3(KEYINPUT64), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G71gat), .B(G78gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT11), .B(new_n509_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n494_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n511_), .A2(new_n512_), .A3(new_n494_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n492_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n511_), .A2(new_n512_), .A3(new_n494_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n517_), .A2(new_n513_), .A3(KEYINPUT72), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n477_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n492_), .A3(new_n515_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT72), .B1(new_n517_), .B2(new_n513_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n468_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n522_), .A3(KEYINPUT74), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G127gat), .B(G155gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G183gat), .B(G211gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n519_), .A2(new_n522_), .A3(KEYINPUT74), .A4(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n491_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n530_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n528_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n519_), .A2(new_n491_), .A3(new_n522_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n541_));
  INV_X1    g340(.A(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(KEYINPUT9), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT6), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(G99gat), .A3(G106gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n546_), .A2(KEYINPUT9), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n544_), .A2(new_n547_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n545_), .A2(new_n546_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n549_), .A2(new_n551_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT7), .ZN(new_n559_));
  INV_X1    g358(.A(G99gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n542_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n557_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT8), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n550_), .B1(G99gat), .B2(G106gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n548_), .A2(KEYINPUT6), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n562_), .B(new_n561_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT8), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n557_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n471_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT34), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n573_), .B(new_n578_), .C1(new_n476_), .C2(new_n571_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n573_), .B1(new_n476_), .B2(new_n571_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n578_), .B(KEYINPUT68), .Z(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n577_), .B2(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT69), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT69), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n583_), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n580_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n591_), .B(KEYINPUT36), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT70), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n593_), .B1(new_n588_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT37), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n593_), .B(new_n598_), .C1(new_n588_), .C2(new_n594_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n540_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT75), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n511_), .A2(new_n512_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n562_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AOI211_X1 g407(.A(KEYINPUT8), .B(new_n556_), .C1(new_n608_), .C2(new_n552_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n569_), .B1(new_n568_), .B2(new_n557_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n554_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n571_), .A2(new_n604_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n603_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT65), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n571_), .B2(new_n604_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT67), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT67), .B(new_n617_), .C1(new_n571_), .C2(new_n604_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n611_), .A2(KEYINPUT12), .A3(new_n512_), .A4(new_n511_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT66), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n605_), .A2(KEYINPUT66), .A3(KEYINPUT12), .A4(new_n611_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n622_), .A2(new_n627_), .A3(new_n603_), .A4(new_n613_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n616_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT5), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n631_), .B(new_n632_), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n616_), .A2(new_n628_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT13), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(KEYINPUT13), .A3(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n490_), .A2(new_n602_), .A3(new_n642_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n643_), .A2(G1gat), .A3(new_n445_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n593_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n458_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n540_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n650_), .A2(new_n489_), .A3(new_n641_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n445_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n644_), .A2(new_n645_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT99), .ZN(G1324gat));
  INV_X1    g455(.A(new_n455_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n643_), .A2(G8gat), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n649_), .A2(new_n455_), .A3(new_n651_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(G8gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n660_), .A3(G8gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n659_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n658_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n664_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n668_), .B2(new_n662_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT39), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n668_), .A2(KEYINPUT101), .A3(new_n662_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n667_), .B(KEYINPUT40), .C1(new_n671_), .C2(new_n670_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  INV_X1    g475(.A(new_n271_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G15gat), .B1(new_n652_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n643_), .A2(G15gat), .A3(new_n677_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT102), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n652_), .B2(new_n451_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n451_), .A2(G22gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n643_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT103), .ZN(G1327gat));
  NAND2_X1  g486(.A1(new_n650_), .A2(new_n648_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT106), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n641_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n490_), .ZN(new_n691_));
  OR3_X1    g490(.A1(new_n691_), .A2(G29gat), .A3(new_n445_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  INV_X1    g493(.A(new_n600_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n694_), .B(new_n695_), .C1(new_n453_), .C2(new_n457_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT104), .ZN(new_n697_));
  INV_X1    g496(.A(new_n456_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n430_), .A2(new_n379_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT98), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n430_), .A2(KEYINPUT98), .A3(new_n379_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n703_), .A3(new_n454_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n454_), .A2(new_n445_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n451_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n703_), .A2(new_n706_), .B1(new_n451_), .B2(new_n450_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n707_), .B2(new_n271_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n694_), .A4(new_n695_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n695_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT43), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n697_), .A2(new_n710_), .A3(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n540_), .A2(new_n641_), .A3(new_n489_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n714_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n693_), .B1(new_n717_), .B2(new_n323_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n714_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n714_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n721_), .A2(new_n693_), .A3(new_n323_), .A4(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G29gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n692_), .B1(new_n718_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT107), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n692_), .C1(new_n718_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1328gat));
  NAND2_X1  g528(.A1(new_n721_), .A2(new_n722_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G36gat), .B1(new_n730_), .B2(new_n657_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n657_), .A2(G36gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n690_), .A2(new_n490_), .A3(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(G1329gat));
  NAND3_X1  g536(.A1(new_n717_), .A2(G43gat), .A3(new_n271_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n691_), .A2(new_n677_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(G43gat), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1330gat));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n717_), .A2(new_n422_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(G50gat), .ZN(new_n745_));
  INV_X1    g544(.A(G50gat), .ZN(new_n746_));
  AOI211_X1 g545(.A(KEYINPUT109), .B(new_n746_), .C1(new_n717_), .C2(new_n422_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n422_), .A2(new_n746_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n745_), .A2(new_n747_), .B1(new_n691_), .B2(new_n748_), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n458_), .A2(new_n488_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n602_), .A3(new_n641_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n497_), .B1(new_n751_), .B2(new_n445_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT110), .Z(new_n753_));
  NAND2_X1  g552(.A1(new_n708_), .A2(new_n647_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n488_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n641_), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n754_), .A2(KEYINPUT111), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT111), .B1(new_n754_), .B2(new_n756_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n445_), .A2(new_n497_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n753_), .B1(new_n759_), .B2(new_n760_), .ZN(G1332gat));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n455_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G64gat), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT48), .B(new_n495_), .C1(new_n759_), .C2(new_n455_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n455_), .A2(new_n495_), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n764_), .A2(new_n765_), .B1(new_n751_), .B2(new_n766_), .ZN(G1333gat));
  OR3_X1    g566(.A1(new_n751_), .A2(G71gat), .A3(new_n677_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n759_), .A2(new_n271_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G71gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G71gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT112), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1334gat));
  OR3_X1    g576(.A1(new_n751_), .A2(G78gat), .A3(new_n451_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n759_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G78gat), .B1(new_n779_), .B2(new_n451_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT50), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1335gat));
  NOR3_X1   g582(.A1(new_n642_), .A2(new_n540_), .A3(new_n488_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n713_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n445_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n689_), .A2(new_n642_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n750_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n445_), .A2(G85gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(G1336gat));
  OAI21_X1  g589(.A(G92gat), .B1(new_n785_), .B2(new_n657_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n657_), .A2(G92gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n788_), .B2(new_n792_), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n785_), .B2(new_n677_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n271_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n788_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n713_), .A2(new_n422_), .A3(new_n784_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n422_), .A2(new_n542_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n800_), .A2(new_n801_), .B1(new_n788_), .B2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g603(.A1(new_n677_), .A2(new_n445_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n657_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n636_), .A2(new_n488_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT114), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n628_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n628_), .A2(KEYINPUT115), .A3(new_n810_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n613_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n603_), .B1(new_n816_), .B2(new_n622_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n813_), .A2(new_n814_), .A3(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n816_), .A2(KEYINPUT55), .A3(new_n603_), .A4(new_n622_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT116), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT56), .B(new_n633_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n622_), .A2(new_n627_), .A3(new_n613_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n603_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n817_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n814_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n633_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n809_), .B1(new_n823_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n472_), .A2(new_n473_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n478_), .A2(new_n479_), .A3(new_n474_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n485_), .A3(new_n834_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n487_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n637_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n832_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n647_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n840_), .B(new_n648_), .C1(new_n832_), .C2(new_n837_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n636_), .A2(new_n836_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n633_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n843_), .B1(new_n846_), .B2(new_n822_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT58), .B1(new_n847_), .B2(KEYINPUT117), .ZN(new_n848_));
  INV_X1    g647(.A(new_n843_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n823_), .B2(new_n831_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n695_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n540_), .B1(new_n842_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n600_), .A2(new_n640_), .A3(new_n639_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n755_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n755_), .A2(new_n857_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n451_), .B(new_n807_), .C1(new_n855_), .C2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n488_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n808_), .B(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n846_), .B2(new_n822_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n837_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n647_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n840_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n647_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n854_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n650_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n863_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n422_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT59), .A3(new_n807_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n489_), .B1(new_n869_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n867_), .B1(new_n882_), .B2(new_n866_), .ZN(G1340gat));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n642_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n865_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n884_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n642_), .B1(new_n869_), .B2(new_n881_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n884_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n865_), .A2(new_n889_), .A3(new_n540_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n650_), .B1(new_n869_), .B2(new_n881_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1342gat));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893_));
  INV_X1    g692(.A(G134gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n600_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n869_), .B2(new_n881_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G134gat), .B1(new_n865_), .B2(new_n648_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n893_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT59), .B1(new_n880_), .B2(new_n807_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n863_), .B1(new_n650_), .B2(new_n877_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n901_), .A2(new_n868_), .A3(new_n422_), .A4(new_n806_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n895_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n894_), .B1(new_n864_), .B2(new_n647_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(KEYINPUT118), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n899_), .A2(new_n905_), .ZN(G1343gat));
  NAND2_X1  g705(.A1(new_n878_), .A2(new_n879_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n271_), .A2(new_n451_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n909_), .A2(new_n455_), .A3(new_n445_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n907_), .A2(KEYINPUT119), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912_));
  INV_X1    g711(.A(new_n910_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n901_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n488_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n641_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT120), .B(G148gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1345gat));
  NAND2_X1  g719(.A1(new_n915_), .A2(new_n540_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1346gat));
  INV_X1    g722(.A(new_n915_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G162gat), .B1(new_n924_), .B2(new_n600_), .ZN(new_n925_));
  INV_X1    g724(.A(G162gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n915_), .A2(new_n926_), .A3(new_n648_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n907_), .A2(new_n451_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n455_), .A2(new_n445_), .A3(new_n271_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n929_), .A2(new_n489_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  XOR2_X1   g731(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n933_));
  NAND3_X1  g732(.A1(new_n932_), .A2(G169gat), .A3(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT121), .A2(KEYINPUT62), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n931_), .B2(new_n219_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n931_), .A2(new_n203_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n934_), .A2(new_n936_), .A3(new_n937_), .ZN(G1348gat));
  NOR2_X1   g737(.A1(new_n929_), .A2(new_n930_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n641_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n353_), .A2(new_n354_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n650_), .A2(new_n930_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n880_), .A2(new_n942_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n451_), .B(new_n944_), .C1(new_n855_), .C2(new_n863_), .ZN(new_n946_));
  AOI21_X1  g745(.A(KEYINPUT122), .B1(new_n946_), .B2(new_n208_), .ZN(new_n947_));
  AND4_X1   g746(.A1(new_n451_), .A2(new_n907_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(KEYINPUT123), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n951_), .B(new_n945_), .C1(new_n947_), .C2(new_n948_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n939_), .A2(new_n351_), .A3(new_n648_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n929_), .A2(new_n600_), .A3(new_n930_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n209_), .ZN(G1351gat));
  NAND3_X1  g755(.A1(new_n455_), .A2(new_n445_), .A3(new_n908_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n901_), .A2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n488_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(KEYINPUT124), .B(G197gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1352gat));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(G204gat), .ZN(new_n963_));
  XOR2_X1   g762(.A(KEYINPUT125), .B(G204gat), .Z(new_n964_));
  NAND2_X1  g763(.A1(new_n958_), .A2(new_n641_), .ZN(new_n965_));
  MUX2_X1   g764(.A(new_n963_), .B(new_n964_), .S(new_n965_), .Z(G1353gat));
  NOR3_X1   g765(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n967_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n958_), .A2(new_n540_), .A3(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(KEYINPUT127), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n969_), .B(new_n971_), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n958_), .A2(new_n337_), .A3(new_n648_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n901_), .A2(new_n600_), .A3(new_n957_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n974_), .B2(new_n337_), .ZN(G1355gat));
endmodule


