//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .A3(new_n202_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(KEYINPUT65), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n217_), .A2(KEYINPUT10), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(KEYINPUT10), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n216_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT6), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n226_), .A2(new_n213_), .A3(KEYINPUT9), .A4(new_n210_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n215_), .A2(new_n220_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n217_), .A2(new_n216_), .A3(KEYINPUT66), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n231_), .A2(new_n217_), .A3(new_n216_), .A4(KEYINPUT66), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n226_), .A2(KEYINPUT67), .A3(new_n210_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n209_), .B(new_n228_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT12), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n228_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n233_), .A2(new_n235_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT8), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n243_), .B1(new_n248_), .B2(new_n209_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n228_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n209_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n243_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n242_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT64), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n248_), .A2(new_n209_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n238_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G120gat), .B(G148gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT5), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(G176gat), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269_));
  INV_X1    g068(.A(new_n267_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n258_), .A2(new_n261_), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n262_), .A2(KEYINPUT69), .A3(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT13), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .A4(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G113gat), .B(G141gat), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G197gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G29gat), .B(G36gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G43gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(G29gat), .A2(G36gat), .ZN(new_n289_));
  INV_X1    g088(.A(G43gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G29gat), .A2(G36gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n288_), .A2(G50gat), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(G50gat), .B1(new_n288_), .B2(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G1gat), .A2(G8gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(KEYINPUT14), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n305_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n295_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n306_), .B(new_n309_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n310_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n288_), .A2(new_n292_), .ZN(new_n318_));
  INV_X1    g117(.A(G50gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n288_), .A2(G50gat), .A3(new_n292_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(KEYINPUT80), .A3(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n314_), .A2(new_n316_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT81), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT15), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(KEYINPUT15), .A3(new_n321_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n317_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n315_), .A3(new_n311_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n324_), .B1(new_n325_), .B2(new_n331_), .ZN(new_n332_));
  AND4_X1   g131(.A1(new_n325_), .A2(new_n314_), .A3(new_n316_), .A4(new_n323_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n286_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n286_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n331_), .A2(new_n325_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n335_), .B(new_n336_), .C1(new_n337_), .C2(new_n324_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n338_), .A3(KEYINPUT82), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(new_n286_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n281_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n345_));
  INV_X1    g144(.A(G211gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT16), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n347_), .B(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(G183gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n346_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n349_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(G211gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n345_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n359_));
  OAI211_X1 g158(.A(G231gat), .B(G233gat), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n357_), .ZN(new_n361_));
  AOI21_X1  g160(.A(G211gat), .B1(new_n355_), .B2(new_n356_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT17), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G231gat), .A2(G233gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT77), .A3(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n360_), .A2(new_n209_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n209_), .B1(new_n360_), .B2(new_n365_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n317_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n363_), .A2(KEYINPUT77), .A3(new_n364_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n364_), .B1(new_n363_), .B2(KEYINPUT77), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n251_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n360_), .A2(new_n365_), .A3(new_n209_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n310_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n354_), .A2(new_n345_), .A3(new_n357_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n344_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT101), .Z(new_n377_));
  XNOR2_X1  g176(.A(G190gat), .B(G218gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n380_), .A2(G134gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(G134gat), .ZN(new_n382_));
  INV_X1    g181(.A(G162gat), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT36), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(KEYINPUT36), .A3(new_n386_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(KEYINPUT74), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G232gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT34), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n329_), .A2(new_n250_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT72), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n250_), .B2(new_n322_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT35), .B(new_n393_), .C1(new_n394_), .C2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT72), .B1(new_n248_), .B2(new_n295_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(KEYINPUT35), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n329_), .A2(new_n250_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n393_), .A2(KEYINPUT35), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n391_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n405_));
  INV_X1    g204(.A(new_n389_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n390_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT73), .B1(new_n403_), .B2(new_n389_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT73), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n406_), .A2(new_n397_), .A3(new_n411_), .A4(new_n402_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G169gat), .A2(G176gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT87), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT22), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G169gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n283_), .A2(KEYINPUT22), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT88), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT88), .B1(new_n283_), .B2(KEYINPUT22), .ZN(new_n421_));
  INV_X1    g220(.A(G176gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n416_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G183gat), .A2(G190gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT23), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT83), .B(G183gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(G190gat), .B2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n416_), .B(KEYINPUT89), .C1(new_n420_), .C2(new_n423_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n426_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT25), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT85), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT25), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G190gat), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n437_), .A2(G183gat), .B1(KEYINPUT26), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT26), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G190gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT84), .B1(new_n429_), .B2(new_n433_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n349_), .A2(KEYINPUT83), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n349_), .A2(KEYINPUT83), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n445_), .B(KEYINPUT25), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n439_), .A2(new_n443_), .A3(new_n444_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n283_), .A2(new_n422_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT24), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n428_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n415_), .A2(KEYINPUT87), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n415_), .A2(KEYINPUT87), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n449_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n432_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n432_), .B2(new_n458_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n461_), .A2(KEYINPUT90), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n432_), .A2(new_n458_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT30), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n467_), .B2(new_n460_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT31), .B1(new_n468_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G127gat), .ZN(new_n476_));
  INV_X1    g275(.A(G134gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G127gat), .A2(G134gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(G113gat), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  INV_X1    g284(.A(G113gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n481_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n484_), .A2(new_n487_), .A3(G120gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(G120gat), .B1(new_n484_), .B2(new_n487_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT90), .B1(new_n461_), .B2(new_n462_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT31), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n473_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n475_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n492_), .B1(new_n475_), .B2(new_n495_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n464_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n475_), .A2(new_n495_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n491_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n475_), .A2(new_n495_), .A3(new_n492_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n463_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G78gat), .B(G106gat), .Z(new_n504_));
  INV_X1    g303(.A(KEYINPUT21), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n285_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(G197gat), .B2(new_n266_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n266_), .A2(G197gat), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n505_), .B(new_n506_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT94), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n285_), .A2(G204gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n285_), .A2(G204gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n507_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G211gat), .B(G218gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT21), .B1(new_n509_), .B2(new_n513_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n514_), .B2(new_n506_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT21), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(G155gat), .A2(G162gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G155gat), .A2(G162gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(G141gat), .A2(G148gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT3), .Z(new_n528_));
  NAND2_X1  g327(.A1(G141gat), .A2(G148gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT2), .Z(new_n530_));
  OAI211_X1 g329(.A(new_n525_), .B(new_n526_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n527_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n526_), .B(KEYINPUT1), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n532_), .B(new_n529_), .C1(new_n533_), .C2(new_n524_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT29), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n523_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G228gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT92), .Z(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n523_), .A2(new_n536_), .A3(new_n539_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n504_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n504_), .A3(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n535_), .A2(KEYINPUT29), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT28), .B(G22gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n319_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n547_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n543_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n544_), .A2(new_n551_), .A3(new_n545_), .A4(new_n550_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n503_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT27), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n523_), .A2(new_n466_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G226gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT19), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n428_), .B1(G183gat), .B2(G190gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n418_), .A2(new_n419_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT98), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n565_), .B(new_n416_), .C1(new_n567_), .C2(G176gat), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n452_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n428_), .A2(new_n451_), .A3(KEYINPUT97), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT25), .B(G183gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n438_), .A2(KEYINPUT26), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n441_), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n453_), .B1(G169gat), .B2(G176gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n568_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(new_n523_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n523_), .A2(new_n466_), .A3(KEYINPUT99), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n561_), .A2(new_n564_), .A3(new_n578_), .A4(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G8gat), .B(G36gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT18), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G64gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(G92gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n563_), .B(KEYINPUT96), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n577_), .A2(new_n523_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT20), .B1(new_n523_), .B2(new_n466_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n580_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n584_), .B1(new_n580_), .B2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n557_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n535_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n484_), .A2(new_n487_), .ZN(new_n593_));
  INV_X1    g392(.A(G120gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n595_), .A2(new_n488_), .A3(new_n534_), .A4(new_n531_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(new_n596_), .A3(KEYINPUT4), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G225gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT4), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n600_), .B(new_n535_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n592_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G1gat), .B(G29gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G85gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT0), .ZN(new_n607_));
  INV_X1    g406(.A(G57gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n602_), .A2(new_n609_), .A3(new_n603_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n580_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n586_), .A2(new_n587_), .A3(new_n585_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n559_), .A2(new_n560_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n617_), .A2(new_n578_), .A3(KEYINPUT20), .A4(new_n579_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n616_), .B1(new_n563_), .B2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT27), .B(new_n615_), .C1(new_n619_), .C2(new_n584_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n591_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n556_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n553_), .A2(new_n554_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n592_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n610_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n612_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n590_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n612_), .A2(new_n630_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .A4(new_n615_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n584_), .A2(KEYINPUT32), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n580_), .A2(new_n635_), .A3(new_n588_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n613_), .B(new_n636_), .C1(new_n635_), .C2(new_n619_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n637_), .A3(new_n555_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n503_), .ZN(new_n639_));
  AND4_X1   g438(.A1(new_n624_), .A2(new_n626_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n503_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n624_), .B1(new_n641_), .B2(new_n638_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n623_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n377_), .A2(new_n414_), .A3(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n614_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT75), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n413_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n414_), .A2(new_n648_), .A3(KEYINPUT37), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n408_), .A2(new_n404_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT75), .B1(new_n410_), .B2(new_n412_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT78), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n375_), .A2(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n368_), .A2(new_n373_), .A3(KEYINPUT78), .A4(new_n374_), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n649_), .A2(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n279_), .A2(new_n280_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT79), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(new_n643_), .A3(new_n342_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n297_), .A3(new_n613_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(KEYINPUT102), .A3(new_n646_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT102), .B1(new_n662_), .B2(new_n646_), .ZN(new_n665_));
  OAI221_X1 g464(.A(new_n645_), .B1(new_n646_), .B2(new_n662_), .C1(new_n664_), .C2(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(new_n644_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n591_), .A2(new_n620_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n298_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n671_), .A3(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n661_), .A2(new_n298_), .A3(new_n669_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G8gat), .B1(new_n644_), .B2(new_n668_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n675_), .A2(KEYINPUT40), .A3(new_n678_), .A4(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(G15gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n661_), .A2(new_n684_), .A3(new_n503_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G15gat), .B1(new_n644_), .B2(new_n639_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT104), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT104), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n687_), .A2(KEYINPUT41), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n687_), .B2(new_n688_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(G1326gat));
  OAI21_X1  g490(.A(G22gat), .B1(new_n644_), .B2(new_n555_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT42), .ZN(new_n693_));
  INV_X1    g492(.A(G22gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n661_), .A2(new_n694_), .A3(new_n625_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n655_), .A2(new_n656_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n414_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n643_), .A2(new_n344_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G29gat), .B1(new_n699_), .B2(new_n613_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n626_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT100), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n641_), .A2(new_n624_), .A3(new_n638_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n622_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n649_), .A2(new_n653_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT105), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT43), .ZN(new_n707_));
  INV_X1    g506(.A(new_n697_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT105), .B(new_n709_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n707_), .A2(new_n708_), .A3(new_n344_), .A4(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(G29gat), .A3(new_n613_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n711_), .A2(new_n712_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n700_), .B1(new_n715_), .B2(new_n716_), .ZN(G1328gat));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n718_), .A3(new_n669_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n668_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n713_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT46), .B(new_n720_), .C1(new_n722_), .C2(new_n718_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n713_), .B2(new_n721_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n720_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1329gat));
  NAND4_X1  g527(.A1(new_n713_), .A2(G43gat), .A3(new_n503_), .A4(new_n716_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n699_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n290_), .B1(new_n730_), .B2(new_n639_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT47), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n734_), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n699_), .B2(new_n625_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n713_), .A2(G50gat), .A3(new_n625_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n739_), .B2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n658_), .A2(new_n342_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n643_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n657_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n613_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n414_), .A3(new_n697_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n746_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1332gat));
  OAI21_X1  g547(.A(G64gat), .B1(new_n746_), .B2(new_n668_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT48), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n668_), .A2(G64gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n743_), .B2(new_n751_), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n746_), .B2(new_n639_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n639_), .A2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n743_), .B2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n746_), .B2(new_n555_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n555_), .A2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n743_), .B2(new_n759_), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n742_), .A2(new_n698_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n613_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n707_), .A2(new_n708_), .A3(new_n710_), .A4(new_n741_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT106), .Z(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(new_n613_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n766_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n762_), .B2(new_n669_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n669_), .A2(G92gat), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT107), .Z(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n765_), .B2(new_n770_), .ZN(G1337gat));
  OAI211_X1 g570(.A(new_n742_), .B(new_n698_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n773_));
  OR3_X1    g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n639_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(new_n639_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G99gat), .B1(new_n764_), .B2(new_n639_), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT109), .B(KEYINPUT51), .C1(new_n776_), .C2(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n779_));
  NAND2_X1  g578(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n780_));
  AND4_X1   g579(.A1(new_n779_), .A2(new_n776_), .A3(new_n780_), .A4(new_n777_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n778_), .A2(new_n781_), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n762_), .A2(new_n216_), .A3(new_n625_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  INV_X1    g583(.A(new_n705_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n643_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n709_), .B1(new_n786_), .B2(KEYINPUT105), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT105), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n788_), .B(KEYINPUT43), .C1(new_n643_), .C2(new_n785_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(new_n708_), .A3(new_n625_), .A4(new_n741_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n784_), .B1(new_n791_), .B2(G106gat), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n784_), .B(G106gat), .C1(new_n764_), .C2(new_n555_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n783_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT53), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n783_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1339gat));
  OAI21_X1  g598(.A(KEYINPUT55), .B1(new_n254_), .B2(new_n257_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n258_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n254_), .A2(KEYINPUT55), .A3(new_n257_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n270_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n267_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n803_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n804_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n314_), .A2(new_n315_), .A3(new_n323_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n286_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT111), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n330_), .A2(new_n316_), .A3(new_n311_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n816_), .A3(new_n286_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n818_), .A2(KEYINPUT112), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(KEYINPUT112), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n271_), .A4(new_n338_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT58), .B1(new_n811_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT115), .B1(new_n823_), .B2(new_n705_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n807_), .A2(new_n805_), .A3(new_n808_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n803_), .B2(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n821_), .B1(new_n827_), .B2(new_n804_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT58), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n785_), .C1(new_n828_), .C2(KEYINPUT58), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  INV_X1    g632(.A(new_n804_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n342_), .B(new_n271_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n819_), .A2(new_n820_), .A3(new_n338_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n837_), .A2(new_n274_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n650_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n833_), .B1(new_n839_), .B2(KEYINPUT113), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n274_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n271_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n807_), .A2(new_n808_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n804_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n845_), .B2(new_n342_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n841_), .B(KEYINPUT57), .C1(new_n846_), .C2(new_n650_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n840_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n832_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n375_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n657_), .A2(new_n658_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .A4(new_n343_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n657_), .A2(new_n658_), .A3(new_n343_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT54), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT110), .B1(new_n856_), .B2(KEYINPUT54), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n851_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n669_), .A2(new_n614_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n556_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n486_), .B1(new_n864_), .B2(new_n343_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n865_), .A2(KEYINPUT116), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(KEYINPUT116), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n849_), .A2(new_n708_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n859_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n863_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT117), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(KEYINPUT59), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n869_), .A2(new_n874_), .A3(new_n870_), .A4(new_n863_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n343_), .A2(new_n486_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n872_), .A2(new_n873_), .A3(new_n875_), .A4(new_n876_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n866_), .A2(new_n867_), .A3(new_n877_), .ZN(G1340gat));
  XOR2_X1   g677(.A(KEYINPUT118), .B(G120gat), .Z(new_n879_));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n658_), .B2(new_n879_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n860_), .A2(new_n863_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n883_), .B2(new_n880_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n872_), .A2(new_n873_), .A3(new_n875_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n658_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(G1341gat));
  OAI21_X1  g687(.A(G127gat), .B1(new_n885_), .B2(new_n850_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n860_), .A2(new_n476_), .A3(new_n697_), .A4(new_n863_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1342gat));
  NAND2_X1  g690(.A1(new_n785_), .A2(G134gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT120), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n477_), .B1(new_n864_), .B2(new_n414_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(KEYINPUT119), .B(new_n477_), .C1(new_n864_), .C2(new_n414_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n886_), .A2(new_n893_), .B1(new_n896_), .B2(new_n897_), .ZN(G1343gat));
  AOI21_X1  g697(.A(new_n555_), .B1(new_n851_), .B2(new_n859_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n639_), .A4(new_n861_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n375_), .B1(new_n832_), .B2(new_n848_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n855_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n625_), .B(new_n639_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT121), .B1(new_n904_), .B2(new_n862_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n343_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(G141gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1344gat));
  AOI21_X1  g707(.A(new_n658_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n909_));
  INV_X1    g708(.A(G148gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1345gat));
  AOI21_X1  g710(.A(new_n708_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT61), .B(G155gat), .Z(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1346gat));
  NAND2_X1  g713(.A1(new_n901_), .A2(new_n905_), .ZN(new_n915_));
  AOI21_X1  g714(.A(G162gat), .B1(new_n915_), .B2(new_n650_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n705_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(G162gat), .B2(new_n917_), .ZN(G1347gat));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n668_), .A2(new_n613_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n556_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n869_), .A2(new_n919_), .A3(new_n342_), .A4(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n697_), .B1(new_n832_), .B2(new_n848_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n342_), .B(new_n922_), .C1(new_n924_), .C2(new_n903_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT122), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n923_), .A2(new_n926_), .A3(G169gat), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n923_), .A2(new_n926_), .A3(KEYINPUT123), .A4(G169gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(KEYINPUT62), .A3(new_n930_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n925_), .A2(new_n567_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n927_), .A2(new_n928_), .A3(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n931_), .A2(new_n932_), .A3(new_n934_), .ZN(G1348gat));
  AND2_X1   g734(.A1(new_n869_), .A2(new_n922_), .ZN(new_n936_));
  AOI21_X1  g735(.A(G176gat), .B1(new_n936_), .B2(new_n281_), .ZN(new_n937_));
  AOI211_X1 g736(.A(new_n422_), .B(new_n658_), .C1(new_n851_), .C2(new_n859_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n922_), .B2(new_n938_), .ZN(G1349gat));
  NOR2_X1   g738(.A1(new_n850_), .A2(new_n572_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n860_), .A2(new_n697_), .A3(new_n922_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n429_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n936_), .A2(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(KEYINPUT124), .ZN(G1350gat));
  AND3_X1   g743(.A1(new_n650_), .A2(new_n441_), .A3(new_n573_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n936_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n869_), .A2(new_n922_), .ZN(new_n947_));
  OAI21_X1  g746(.A(G190gat), .B1(new_n947_), .B2(new_n705_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1351gat));
  NOR2_X1   g750(.A1(new_n904_), .A2(new_n921_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n342_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n281_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n899_), .A2(new_n375_), .A3(new_n639_), .A4(new_n920_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n959_), .A2(KEYINPUT126), .A3(new_n961_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n904_), .A2(new_n850_), .A3(new_n921_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n960_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n958_), .B1(new_n962_), .B2(new_n965_), .ZN(new_n966_));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n959_), .B2(new_n961_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n964_), .A2(new_n963_), .A3(new_n960_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n967_), .A2(new_n957_), .A3(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n966_), .A2(new_n969_), .ZN(G1354gat));
  NAND3_X1  g769(.A1(new_n952_), .A2(G218gat), .A3(new_n785_), .ZN(new_n971_));
  NOR3_X1   g770(.A1(new_n904_), .A2(new_n414_), .A3(new_n921_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n971_), .B1(new_n972_), .B2(G218gat), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n971_), .B(KEYINPUT127), .C1(new_n972_), .C2(G218gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(G1355gat));
endmodule


