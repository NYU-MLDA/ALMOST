//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G106gat), .Z(new_n213_));
  AOI22_X1  g012(.A1(new_n212_), .A2(new_n213_), .B1(new_n202_), .B2(KEYINPUT9), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT9), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n208_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n202_), .A2(KEYINPUT8), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n208_), .B1(new_n205_), .B2(KEYINPUT65), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n203_), .B(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n221_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(KEYINPUT12), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G230gat), .A2(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G120gat), .B(G148gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT5), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G176gat), .B(G204gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n235_), .A2(new_n237_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n242_), .B(new_n247_), .C1(new_n241_), .C2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n241_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n241_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n246_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT13), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(KEYINPUT13), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT66), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT35), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G29gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT68), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G43gat), .B(G50gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n267_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n269_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n227_), .A2(new_n276_), .B1(new_n264_), .B2(new_n263_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n266_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n275_), .B(KEYINPUT15), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n277_), .B1(new_n280_), .B2(new_n227_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  OAI221_X1 g081(.A(new_n277_), .B1(new_n278_), .B2(new_n266_), .C1(new_n280_), .C2(new_n227_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n287_), .B(KEYINPUT36), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n284_), .A2(KEYINPUT71), .A3(new_n290_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n289_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT37), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n289_), .A2(new_n297_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n296_), .A2(new_n297_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n234_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT72), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  OR2_X1    g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT17), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n302_), .A2(new_n309_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G127gat), .B(G155gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT16), .ZN(new_n314_));
  XOR2_X1   g113(.A(G183gat), .B(G211gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .A4(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT73), .B1(new_n310_), .B2(new_n312_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n316_), .A2(new_n311_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  AOI211_X1 g120(.A(KEYINPUT73), .B(new_n321_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n317_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n299_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT95), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT19), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT77), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(G169gat), .B2(G176gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT78), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT78), .B1(new_n339_), .B2(new_n341_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n336_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n336_), .B1(G169gat), .B2(G176gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n342_), .A3(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT75), .B(G183gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(KEYINPUT76), .A2(G190gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT26), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT23), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n345_), .A2(new_n350_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G169gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n359_), .ZN(new_n363_));
  INV_X1    g162(.A(G190gat), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n352_), .A2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n362_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT21), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(G197gat), .B2(G204gat), .ZN(new_n369_));
  OR2_X1    g168(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(new_n372_), .B2(G204gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n372_), .B2(G204gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n373_), .B(new_n374_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n368_), .B1(new_n374_), .B2(KEYINPUT90), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n376_), .B(new_n379_), .C1(KEYINPUT90), .C2(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n335_), .B1(new_n367_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(KEYINPUT91), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n359_), .B1(G183gat), .B2(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n362_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n346_), .A2(new_n336_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n350_), .A2(new_n359_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n378_), .A2(new_n380_), .A3(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n383_), .A2(new_n385_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n334_), .B1(new_n382_), .B2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n378_), .A2(new_n380_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(KEYINPUT93), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n350_), .A2(new_n397_), .A3(new_n359_), .A4(new_n388_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n396_), .A2(new_n398_), .B1(new_n362_), .B2(new_n384_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT20), .B(new_n395_), .C1(new_n399_), .C2(new_n394_), .ZN(new_n400_));
  OAI22_X1  g199(.A1(new_n393_), .A2(KEYINPUT99), .B1(new_n400_), .B2(new_n333_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT99), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n402_), .B(new_n334_), .C1(new_n382_), .C2(new_n392_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n331_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  AOI211_X1 g204(.A(new_n335_), .B(new_n333_), .C1(new_n367_), .C2(new_n381_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n394_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n400_), .A2(new_n333_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n408_), .B2(new_n330_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n414_));
  OR2_X1    g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT82), .B1(new_n413_), .B2(KEYINPUT1), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT83), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n413_), .A2(KEYINPUT1), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(KEYINPUT1), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n415_), .A4(new_n414_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G141gat), .B(G148gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT2), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n429_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n415_), .A2(new_n413_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n427_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G127gat), .B(G134gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT81), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G113gat), .B(G120gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n412_), .B1(new_n437_), .B2(new_n441_), .ZN(new_n442_));
  AOI221_X4 g241(.A(KEYINPUT85), .B1(new_n434_), .B2(new_n435_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n427_), .B2(new_n436_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n446_), .B2(new_n441_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n440_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n439_), .B(new_n448_), .ZN(new_n449_));
  NOR4_X1   g248(.A1(new_n443_), .A2(new_n445_), .A3(new_n412_), .A4(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n411_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT0), .B(G57gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n437_), .A2(KEYINPUT85), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n425_), .A2(new_n426_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n444_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n459_), .A3(new_n441_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT96), .B1(new_n449_), .B2(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n457_), .A2(KEYINPUT96), .A3(new_n459_), .A4(new_n441_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n456_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n457_), .A2(new_n456_), .A3(new_n459_), .A4(new_n441_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n411_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n451_), .B(new_n455_), .C1(new_n464_), .C2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n455_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n443_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n463_), .B1(new_n470_), .B2(new_n442_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n471_), .B2(KEYINPUT4), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n466_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n396_), .A2(new_n398_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n394_), .B1(new_n475_), .B2(new_n385_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n395_), .A2(KEYINPUT20), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n333_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n406_), .A2(new_n407_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n330_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n330_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n405_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n410_), .A2(new_n468_), .A3(new_n474_), .A4(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G99gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G43gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n449_), .A2(KEYINPUT31), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n449_), .A2(KEYINPUT31), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G227gat), .A2(G233gat), .ZN(new_n491_));
  INV_X1    g290(.A(G15gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n360_), .B2(new_n366_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n360_), .A2(new_n366_), .A3(new_n494_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n498_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n490_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n490_), .B1(new_n502_), .B2(new_n499_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n486_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n499_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n490_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n485_), .A3(new_n503_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n457_), .A2(KEYINPUT29), .A3(new_n459_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT87), .B(G233gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT86), .B(G228gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n394_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n391_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n390_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n517_), .A2(new_n518_), .B1(new_n458_), .B2(new_n519_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n512_), .A2(new_n516_), .B1(new_n520_), .B2(new_n515_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G78gat), .B(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT28), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n519_), .B(new_n527_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n521_), .A2(new_n523_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n525_), .A2(new_n532_), .A3(KEYINPUT92), .A4(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT92), .B1(new_n521_), .B2(new_n523_), .ZN(new_n536_));
  OAI22_X1  g335(.A1(new_n535_), .A2(new_n524_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n511_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n483_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n471_), .A2(KEYINPUT4), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(KEYINPUT98), .A3(new_n411_), .A4(new_n465_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n465_), .A2(new_n411_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n464_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n455_), .B1(new_n471_), .B2(new_n466_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n468_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n480_), .A2(new_n481_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n467_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n540_), .A2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n455_), .A2(KEYINPUT33), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n451_), .A3(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n546_), .A2(new_n548_), .A3(new_n549_), .A4(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n534_), .A2(new_n537_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n478_), .A2(new_n479_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n400_), .A2(new_n333_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n382_), .A2(new_n392_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n402_), .B1(new_n560_), .B2(new_n334_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n393_), .A2(KEYINPUT99), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n558_), .B1(new_n563_), .B2(new_n557_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n455_), .B1(new_n551_), .B2(new_n451_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n472_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n554_), .A2(new_n555_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n534_), .A2(new_n537_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n511_), .B1(new_n483_), .B2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n539_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n309_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(new_n275_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT74), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n574_), .B(new_n576_), .C1(new_n280_), .C2(new_n309_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n275_), .B(new_n309_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(new_n575_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n576_), .B1(new_n572_), .B2(new_n275_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT15), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n275_), .B(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n587_), .B2(new_n572_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n578_), .A2(new_n575_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n584_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  NOR4_X1   g390(.A1(new_n260_), .A2(new_n324_), .A3(new_n571_), .A4(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n565_), .A2(new_n566_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n304_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT100), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n568_), .A2(new_n570_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n539_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n258_), .A2(new_n591_), .ZN(new_n602_));
  AND4_X1   g401(.A1(new_n601_), .A2(new_n296_), .A3(new_n323_), .A4(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n304_), .B1(new_n603_), .B2(new_n594_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(G1324gat));
  NAND2_X1  g405(.A1(new_n410_), .A2(new_n482_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n592_), .A2(new_n305_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(G8gat), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1325gat));
  AOI21_X1  g414(.A(new_n492_), .B1(new_n603_), .B2(new_n511_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT41), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n592_), .A2(new_n492_), .A3(new_n511_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1326gat));
  INV_X1    g418(.A(G22gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n603_), .B2(new_n569_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n592_), .A2(new_n620_), .A3(new_n569_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(new_n323_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n295_), .ZN(new_n627_));
  NOR4_X1   g426(.A1(new_n571_), .A2(new_n627_), .A3(new_n591_), .A4(new_n258_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n594_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n298_), .A2(new_n291_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n295_), .B2(KEYINPUT37), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT102), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n601_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n571_), .B2(new_n299_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  AND4_X1   g438(.A1(KEYINPUT44), .A2(new_n639_), .A3(new_n626_), .A4(new_n602_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n602_), .A2(new_n626_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT44), .B1(new_n639_), .B2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n594_), .A2(G29gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n629_), .B1(new_n644_), .B2(new_n645_), .ZN(G1328gat));
  INV_X1    g445(.A(G36gat), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n607_), .A2(KEYINPUT103), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n607_), .A2(KEYINPUT103), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n628_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT45), .ZN(new_n652_));
  INV_X1    g451(.A(new_n607_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n640_), .A2(new_n653_), .A3(new_n643_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(new_n647_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n652_), .B(KEYINPUT46), .C1(new_n654_), .C2(new_n647_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1329gat));
  AOI21_X1  g458(.A(G43gat), .B1(new_n628_), .B2(new_n511_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n511_), .A2(G43gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n644_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT47), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1330gat));
  INV_X1    g463(.A(G50gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n628_), .A2(new_n665_), .A3(new_n569_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n640_), .A2(new_n555_), .A3(new_n643_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT104), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n670_), .B(new_n666_), .C1(new_n667_), .C2(new_n665_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1331gat));
  AND2_X1   g471(.A1(new_n256_), .A2(new_n257_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n324_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n583_), .A2(new_n590_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n571_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n678_), .A2(G57gat), .A3(new_n593_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n571_), .A2(new_n295_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(new_n591_), .A3(new_n260_), .A4(new_n323_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n593_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT105), .Z(G1332gat));
  INV_X1    g483(.A(new_n650_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G64gat), .B1(new_n681_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n685_), .A2(G64gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n678_), .B2(new_n689_), .ZN(G1333gat));
  INV_X1    g489(.A(new_n511_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G71gat), .B1(new_n681_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n691_), .A2(G71gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n678_), .B2(new_n695_), .ZN(G1334gat));
  OR3_X1    g495(.A1(new_n678_), .A2(G78gat), .A3(new_n555_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n681_), .A2(new_n555_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(G78gat), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G78gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(G1335gat));
  NOR3_X1   g503(.A1(new_n673_), .A2(new_n323_), .A3(new_n675_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G85gat), .B1(new_n708_), .B2(new_n593_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n676_), .A2(new_n260_), .A3(new_n295_), .A4(new_n626_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n215_), .A3(new_n594_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1336gat));
  OAI21_X1  g512(.A(G92gat), .B1(new_n708_), .B2(new_n685_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n216_), .A3(new_n607_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1337gat));
  OAI21_X1  g515(.A(G99gat), .B1(new_n708_), .B2(new_n691_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n511_), .A2(new_n212_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n710_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n569_), .A3(new_n213_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  INV_X1    g521(.A(G106gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(new_n555_), .B(new_n706_), .C1(new_n635_), .C2(new_n638_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n707_), .B2(new_n569_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n722_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n636_), .B1(new_n601_), .B2(new_n631_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n571_), .A2(new_n299_), .A3(new_n633_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n569_), .B(new_n705_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G106gat), .B1(new_n732_), .B2(KEYINPUT110), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n733_), .A2(KEYINPUT52), .A3(new_n727_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n721_), .B1(new_n729_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n721_), .C1(new_n729_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  NAND3_X1  g538(.A1(new_n238_), .A2(new_n239_), .A3(new_n251_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n242_), .A2(KEYINPUT55), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n247_), .B1(new_n252_), .B2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(KEYINPUT56), .A3(new_n743_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n588_), .A2(new_n589_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n578_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n582_), .B1(new_n750_), .B2(new_n576_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n573_), .A2(new_n576_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n280_), .B2(new_n309_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n749_), .A2(new_n582_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n249_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(KEYINPUT112), .B2(new_n744_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT113), .B1(new_n748_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n631_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT113), .B(KEYINPUT58), .C1(new_n748_), .C2(new_n756_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n254_), .A2(new_n754_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n250_), .A2(new_n252_), .A3(new_n246_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n591_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n249_), .B2(new_n675_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n745_), .A2(new_n747_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n764_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n762_), .B1(new_n771_), .B2(new_n295_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n747_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n744_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n766_), .B1(new_n591_), .B2(new_n765_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n249_), .A2(new_n675_), .A3(KEYINPUT111), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n763_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(KEYINPUT57), .A3(new_n296_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n626_), .B1(new_n761_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n673_), .A2(new_n323_), .A3(new_n591_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n631_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n569_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n593_), .A2(new_n607_), .A3(new_n691_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT115), .B(G113gat), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n591_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n788_), .B2(new_n591_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT114), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n796_), .C1(new_n788_), .C2(new_n591_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n793_), .A2(new_n795_), .B1(new_n798_), .B2(new_n800_), .ZN(G1340gat));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n673_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n789_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n259_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n802_), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n789_), .A2(new_n807_), .A3(new_n323_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n626_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n807_), .ZN(G1342gat));
  AOI21_X1  g609(.A(G134gat), .B1(new_n789_), .B2(new_n295_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT116), .B(G134gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n299_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n793_), .B2(new_n813_), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n781_), .A2(new_n785_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n555_), .A2(new_n511_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n650_), .A2(new_n593_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n591_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n259_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT117), .B(G148gat), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n821_), .B(new_n822_), .Z(G1345gat));
  AOI211_X1 g622(.A(new_n555_), .B(new_n511_), .C1(new_n781_), .C2(new_n785_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n824_), .A2(new_n323_), .A3(new_n817_), .A4(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n818_), .B2(new_n626_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1346gat));
  NOR2_X1   g631(.A1(new_n818_), .A2(new_n299_), .ZN(new_n833_));
  INV_X1    g632(.A(G162gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n295_), .A2(new_n834_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(new_n833_), .A2(new_n834_), .B1(new_n818_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT120), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  OAI221_X1 g637(.A(new_n838_), .B1(new_n818_), .B2(new_n835_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1347gat));
  NAND2_X1  g639(.A1(new_n650_), .A2(new_n593_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n691_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n815_), .A2(new_n675_), .A3(new_n555_), .A4(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT22), .B(G169gat), .Z(new_n844_));
  OR2_X1    g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n337_), .B1(new_n843_), .B2(KEYINPUT121), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n786_), .A2(new_n848_), .A3(new_n675_), .A4(new_n842_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n846_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n845_), .B1(new_n850_), .B2(new_n851_), .ZN(G1348gat));
  OR2_X1    g651(.A1(new_n786_), .A2(KEYINPUT122), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n786_), .A2(KEYINPUT122), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n259_), .A2(new_n338_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n853_), .A2(new_n842_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n815_), .A2(new_n555_), .A3(new_n842_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n338_), .B1(new_n857_), .B2(new_n673_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n856_), .A2(new_n858_), .ZN(G1349gat));
  OR2_X1    g658(.A1(new_n626_), .A2(new_n386_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n857_), .A2(KEYINPUT123), .A3(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT123), .B1(new_n857_), .B2(new_n860_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n853_), .A2(new_n854_), .A3(new_n323_), .A4(new_n842_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n352_), .B2(new_n864_), .ZN(G1350gat));
  OAI21_X1  g664(.A(G190gat), .B1(new_n857_), .B2(new_n299_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n295_), .A2(new_n387_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n857_), .B2(new_n867_), .ZN(G1351gat));
  INV_X1    g667(.A(new_n841_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n824_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n591_), .ZN(new_n871_));
  INV_X1    g670(.A(G197gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1352gat));
  NOR2_X1   g672(.A1(new_n870_), .A2(new_n259_), .ZN(new_n874_));
  INV_X1    g673(.A(G204gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1353gat));
  AOI21_X1  g675(.A(new_n626_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT124), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n870_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1354gat));
  INV_X1    g680(.A(new_n870_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n295_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT125), .B(G218gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n299_), .A2(new_n884_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT126), .Z(new_n886_));
  AOI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n882_), .B2(new_n886_), .ZN(G1355gat));
endmodule


