//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(new_n203_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT76), .B(G176gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G169gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n208_), .A2(new_n209_), .B1(G169gat), .B2(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(new_n205_), .B2(new_n203_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n214_), .A2(new_n218_), .A3(new_n220_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT30), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G71gat), .B(G99gat), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n225_), .B(KEYINPUT30), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G227gat), .A2(G233gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT77), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT78), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n202_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n230_), .A2(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n235_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n202_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n236_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G113gat), .B(G120gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT80), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT31), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(KEYINPUT79), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n239_), .A2(new_n244_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255_));
  XOR2_X1   g054(.A(G155gat), .B(G162gat), .Z(new_n256_));
  INV_X1    g055(.A(G141gat), .ZN(new_n257_));
  INV_X1    g056(.A(G148gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT3), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(KEYINPUT81), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n261_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n256_), .B1(new_n260_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT1), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n256_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n268_), .A2(new_n262_), .A3(new_n259_), .A4(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n266_), .A2(KEYINPUT82), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT82), .B1(new_n266_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n248_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n270_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n247_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT93), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n271_), .A2(new_n272_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n248_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT92), .B1(new_n277_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n273_), .A2(new_n289_), .A3(KEYINPUT4), .A4(new_n276_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n281_), .B1(new_n291_), .B2(new_n280_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G29gat), .ZN(new_n293_));
  INV_X1    g092(.A(G85gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G57gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n255_), .B1(new_n292_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G92gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT18), .B(G64gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n210_), .B1(new_n213_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n215_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT89), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n206_), .B1(new_n311_), .B2(new_n217_), .ZN(new_n312_));
  OR2_X1    g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n223_), .B1(new_n313_), .B2(new_n309_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n308_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G197gat), .B(G204gat), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT21), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT86), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n316_), .A2(KEYINPUT21), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n315_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT19), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n323_), .B2(new_n225_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(KEYINPUT20), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n326_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n315_), .B2(new_n323_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n323_), .A2(new_n225_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n306_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(KEYINPUT91), .B(new_n306_), .C1(new_n329_), .C2(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n333_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n326_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n305_), .A3(new_n328_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT90), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT90), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n340_), .A2(new_n343_), .A3(new_n305_), .A4(new_n328_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n337_), .A2(new_n338_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n291_), .A2(new_n280_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n277_), .B(KEYINPUT96), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n279_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n297_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n299_), .A2(new_n300_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n301_), .A2(new_n345_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n292_), .A2(new_n298_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n292_), .A2(new_n298_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n324_), .A2(KEYINPUT20), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT97), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n323_), .A2(new_n225_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n355_), .A2(new_n356_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n326_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n332_), .A2(new_n333_), .A3(new_n330_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT32), .A3(new_n305_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n340_), .A2(new_n328_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n354_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n254_), .B1(new_n351_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G22gat), .B(G50gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n323_), .B1(new_n372_), .B2(new_n275_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT85), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  OR3_X1    g175(.A1(new_n282_), .A2(KEYINPUT84), .A3(new_n372_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT84), .B1(new_n282_), .B2(new_n372_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n323_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(new_n375_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G78gat), .B(G106gat), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n282_), .A2(new_n383_), .A3(new_n372_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n282_), .B2(new_n372_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n382_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n380_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n380_), .A2(new_n390_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n371_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n371_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n395_), .A2(new_n391_), .A3(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n354_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n397_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n395_), .B2(new_n391_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n254_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n239_), .A2(new_n244_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n250_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n251_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n397_), .B2(new_n394_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT27), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n345_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n341_), .B(KEYINPUT98), .Z(new_n410_));
  AOI21_X1  g209(.A(new_n305_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT27), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n402_), .A2(new_n407_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n368_), .A2(new_n398_), .B1(new_n399_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G190gat), .B(G218gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G134gat), .B(G162gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT36), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G29gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G43gat), .B(G50gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n423_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT64), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT9), .ZN(new_n429_));
  OR2_X1    g228(.A1(G85gat), .A2(G92gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT9), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(KEYINPUT64), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G106gat), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(KEYINPUT10), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(KEYINPUT10), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n439_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n433_), .A2(new_n438_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n440_), .A3(new_n439_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n446_), .A2(new_n436_), .A3(new_n437_), .A4(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT8), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(KEYINPUT65), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n430_), .A2(new_n427_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n444_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n426_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT69), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G232gat), .A2(G233gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT34), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n461_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n448_), .A2(new_n452_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n450_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n444_), .A3(new_n423_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n457_), .A2(new_n463_), .A3(new_n464_), .A4(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT69), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n426_), .B2(new_n455_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n464_), .B(new_n469_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n462_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n420_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n470_), .A2(new_n475_), .A3(KEYINPUT70), .A4(new_n419_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(KEYINPUT36), .A3(new_n418_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n414_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(G57gat), .A2(G64gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G57gat), .A2(G64gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n488_));
  INV_X1    g287(.A(G71gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G78gat), .ZN(new_n490_));
  INV_X1    g289(.A(G78gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G71gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n487_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n488_), .B1(new_n487_), .B2(new_n493_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n485_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(G57gat), .A2(G64gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G57gat), .A2(G64gat), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT11), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G71gat), .B(G78gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT66), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n487_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n496_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G231gat), .A2(G233gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT73), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n506_), .B(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G15gat), .B(G22gat), .Z(new_n510_));
  NAND2_X1  g309(.A1(G1gat), .A2(G8gat), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(KEYINPUT14), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n511_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G1gat), .A2(G8gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n513_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n517_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n509_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G127gat), .B(G155gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G211gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT16), .B(G183gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n523_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n529_), .B2(new_n523_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n468_), .B(new_n444_), .C1(new_n498_), .C2(new_n505_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n503_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n497_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n455_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n536_), .A3(KEYINPUT12), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT12), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n506_), .A2(new_n538_), .A3(new_n455_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G120gat), .B(G148gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT5), .B(G176gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(KEYINPUT67), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n546_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n552_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(KEYINPUT13), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(KEYINPUT13), .B1(new_n553_), .B2(new_n554_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n423_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n520_), .A2(new_n521_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n512_), .B(new_n513_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n517_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n423_), .B1(new_n563_), .B2(new_n519_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n424_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n423_), .A2(new_n424_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G169gat), .B(G197gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(new_n575_), .A3(new_n571_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n558_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n483_), .A2(new_n532_), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n582_), .B2(new_n399_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT99), .ZN(new_n584_));
  INV_X1    g383(.A(new_n367_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n345_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n349_), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n255_), .B(KEYINPUT33), .C1(new_n292_), .C2(new_n298_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n406_), .B(new_n398_), .C1(new_n585_), .C2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n412_), .A2(new_n409_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n407_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n406_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n399_), .B(new_n591_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n482_), .A2(KEYINPUT71), .A3(KEYINPUT37), .ZN(new_n596_));
  OR2_X1    g395(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n597_));
  NAND2_X1  g396(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n480_), .A2(new_n481_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n596_), .A2(new_n532_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n579_), .B(KEYINPUT74), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n558_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(G1gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n354_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT38), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(KEYINPUT38), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n584_), .B(new_n611_), .C1(new_n609_), .C2(new_n607_), .ZN(G1324gat));
  INV_X1    g411(.A(G8gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n591_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n605_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n483_), .A2(new_n532_), .A3(new_n614_), .A4(new_n581_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n616_), .A2(new_n617_), .A3(G8gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n616_), .B2(G8gat), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1325gat));
  INV_X1    g421(.A(G15gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n605_), .A2(new_n623_), .A3(new_n254_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n483_), .A2(new_n532_), .A3(new_n254_), .A4(new_n581_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G15gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT101), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT41), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n629_), .A3(G15gat), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n627_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n628_), .B1(new_n627_), .B2(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n624_), .B1(new_n631_), .B2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n398_), .B(KEYINPUT102), .Z(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n605_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n582_), .B2(new_n635_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT103), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n641_), .B(G22gat), .C1(new_n582_), .C2(new_n635_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n640_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n637_), .B1(new_n643_), .B2(new_n644_), .ZN(G1327gat));
  INV_X1    g444(.A(new_n532_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n595_), .A2(new_n646_), .A3(new_n482_), .A4(new_n604_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT105), .ZN(new_n648_));
  INV_X1    g447(.A(new_n482_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n590_), .B2(new_n594_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n646_), .A4(new_n604_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n354_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n581_), .A2(new_n646_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n596_), .A2(new_n599_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(KEYINPUT104), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n595_), .B2(new_n658_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n658_), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n662_), .B(new_n659_), .C1(new_n590_), .C2(new_n594_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n656_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(G29gat), .A3(new_n354_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n656_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n654_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  OAI21_X1  g468(.A(new_n659_), .B1(new_n414_), .B2(new_n662_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n595_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n655_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n614_), .B1(new_n672_), .B2(KEYINPUT44), .ZN(new_n673_));
  INV_X1    g472(.A(new_n668_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G36gat), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n591_), .A2(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n648_), .A2(new_n652_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n648_), .A2(KEYINPUT45), .A3(new_n652_), .A4(new_n676_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n675_), .A2(KEYINPUT46), .A3(new_n679_), .A4(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n591_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(new_n668_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n680_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(new_n687_), .ZN(G1329gat));
  NAND4_X1  g487(.A1(new_n666_), .A2(new_n668_), .A3(G43gat), .A4(new_n254_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n648_), .A2(new_n254_), .A3(new_n652_), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT47), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(new_n695_), .A3(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1330gat));
  INV_X1    g496(.A(new_n398_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n666_), .A2(new_n668_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G50gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n635_), .A2(G50gat), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT106), .Z(new_n702_));
  NAND2_X1  g501(.A1(new_n653_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1331gat));
  NOR2_X1   g503(.A1(new_n557_), .A2(new_n646_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n483_), .A2(new_n603_), .A3(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT107), .B(G57gat), .Z(new_n707_));
  NOR3_X1   g506(.A1(new_n706_), .A2(new_n399_), .A3(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT108), .Z(new_n709_));
  NAND2_X1  g508(.A1(new_n558_), .A2(new_n580_), .ZN(new_n710_));
  NOR4_X1   g509(.A1(new_n414_), .A2(new_n646_), .A3(new_n658_), .A4(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n354_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n714_), .A3(new_n614_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n483_), .A2(new_n614_), .A3(new_n603_), .A4(new_n705_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT48), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G64gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1333gat));
  NAND3_X1  g521(.A1(new_n711_), .A2(new_n489_), .A3(new_n254_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G71gat), .B1(new_n706_), .B2(new_n406_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(G1334gat));
  NAND3_X1  g526(.A1(new_n711_), .A2(new_n491_), .A3(new_n636_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G78gat), .B1(new_n706_), .B2(new_n635_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT110), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(G78gat), .C1(new_n706_), .C2(new_n635_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n730_), .A2(new_n731_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n731_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n728_), .B1(new_n734_), .B2(new_n735_), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n710_), .A2(new_n532_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n650_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n354_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n737_), .B(KEYINPUT111), .Z(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n399_), .A2(new_n294_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n738_), .B2(new_n614_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n614_), .A2(G92gat), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT112), .Z(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  AOI21_X1  g547(.A(new_n440_), .B1(new_n742_), .B2(new_n254_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n441_), .A2(new_n442_), .ZN(new_n750_));
  AND4_X1   g549(.A1(new_n254_), .A2(new_n650_), .A3(new_n750_), .A4(new_n737_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n753_), .B(new_n754_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n738_), .A2(new_n439_), .A3(new_n698_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n698_), .B(new_n740_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G106gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G106gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n600_), .A2(new_n770_), .A3(new_n557_), .A4(new_n603_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n596_), .A2(new_n557_), .A3(new_n532_), .A4(new_n599_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT54), .B1(new_n772_), .B2(new_n602_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n542_), .A2(new_n545_), .A3(new_n551_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n537_), .A2(new_n544_), .A3(new_n539_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n537_), .A2(KEYINPUT114), .A3(new_n544_), .A4(new_n539_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n542_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n540_), .A2(KEYINPUT55), .A3(new_n541_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT55), .B1(new_n540_), .B2(new_n541_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n782_), .B(new_n544_), .C1(new_n537_), .C2(new_n539_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT115), .A3(new_n781_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n787_), .A2(new_n550_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n550_), .A4(new_n791_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n776_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n559_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n563_), .A2(new_n519_), .A3(new_n423_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n425_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT116), .B1(new_n799_), .B2(new_n566_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n565_), .A2(new_n801_), .A3(new_n567_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n802_), .A3(new_n570_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n560_), .A2(new_n564_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n576_), .B1(new_n804_), .B2(new_n568_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n803_), .A2(KEYINPUT117), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n803_), .B2(new_n805_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n577_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n796_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT58), .B1(new_n796_), .B2(new_n809_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n579_), .A2(new_n775_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n553_), .A2(new_n554_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n803_), .A2(new_n805_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n803_), .A2(KEYINPUT117), .A3(new_n805_), .ZN(new_n819_));
  AND4_X1   g618(.A1(new_n815_), .A2(new_n818_), .A3(new_n577_), .A4(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n649_), .B1(new_n814_), .B2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n649_), .B(new_n822_), .C1(new_n814_), .C2(new_n820_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n812_), .A2(new_n658_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n774_), .B1(new_n826_), .B2(new_n532_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n614_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G113gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT120), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n831_), .A2(KEYINPUT120), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n603_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  AND4_X1   g633(.A1(KEYINPUT115), .A2(new_n781_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT115), .B1(new_n790_), .B2(new_n781_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n837_), .B2(new_n550_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n795_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n809_), .B(new_n775_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n796_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n658_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n813_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n809_), .A2(new_n815_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n822_), .B1(new_n848_), .B2(new_n649_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n825_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n844_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT119), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n824_), .A2(new_n825_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n844_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n646_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n774_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(new_n829_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n830_), .B(new_n834_), .C1(new_n858_), .C2(new_n828_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G113gat), .B1(new_n858_), .B2(new_n579_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1340gat));
  OAI211_X1 g661(.A(new_n558_), .B(new_n830_), .C1(new_n858_), .C2(new_n828_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  AOI21_X1  g664(.A(G120gat), .B1(new_n558_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT121), .B1(new_n865_), .B2(G120gat), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n858_), .B(new_n868_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n864_), .A2(new_n870_), .ZN(G1341gat));
  AND2_X1   g670(.A1(new_n532_), .A2(G127gat), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n830_), .B(new_n872_), .C1(new_n858_), .C2(new_n828_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G127gat), .B1(new_n858_), .B2(new_n532_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1342gat));
  AND2_X1   g675(.A1(new_n658_), .A2(G134gat), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n830_), .B(new_n877_), .C1(new_n858_), .C2(new_n828_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G134gat), .B1(new_n858_), .B2(new_n482_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n614_), .A2(new_n399_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n857_), .A2(new_n592_), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n580_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n257_), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n557_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n258_), .ZN(G1345gat));
  AND2_X1   g686(.A1(new_n771_), .A2(new_n773_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(new_n532_), .A3(new_n592_), .A4(new_n882_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT122), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  INV_X1    g691(.A(G162gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n883_), .A2(new_n893_), .A3(new_n662_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n857_), .A2(new_n592_), .A3(new_n482_), .A4(new_n882_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n893_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(KEYINPUT123), .A3(new_n893_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n894_), .B1(new_n898_), .B2(new_n899_), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n591_), .A2(new_n354_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n406_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n532_), .B1(new_n853_), .B2(new_n844_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n635_), .B(new_n903_), .C1(new_n904_), .C2(new_n888_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905_), .B2(new_n580_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT62), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n579_), .A2(new_n209_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT124), .Z(new_n909_));
  OAI21_X1  g708(.A(new_n907_), .B1(new_n905_), .B2(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(new_n902_), .B1(new_n856_), .B2(new_n774_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n911_), .A2(G176gat), .A3(new_n593_), .A4(new_n558_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n914_));
  INV_X1    g713(.A(new_n905_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n558_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n916_), .A2(new_n208_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n913_), .A2(new_n914_), .A3(new_n917_), .ZN(G1349gat));
  AOI211_X1 g717(.A(new_n402_), .B(new_n902_), .C1(new_n856_), .C2(new_n774_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n919_), .B2(new_n532_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n221_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n827_), .A2(new_n921_), .A3(new_n635_), .A4(new_n903_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT126), .B1(new_n922_), .B2(new_n646_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n915_), .A2(new_n924_), .A3(new_n532_), .A4(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT127), .B1(new_n920_), .B2(new_n926_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n857_), .A2(new_n532_), .A3(new_n593_), .A4(new_n901_), .ZN(new_n928_));
  INV_X1    g727(.A(G183gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n923_), .A4(new_n925_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n927_), .A2(new_n932_), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n905_), .B2(new_n662_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n482_), .A2(new_n222_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n905_), .B2(new_n935_), .ZN(G1351gat));
  NAND3_X1  g735(.A1(new_n911_), .A2(new_n592_), .A3(new_n579_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g737(.A1(new_n911_), .A2(new_n592_), .A3(new_n558_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n911_), .A2(new_n532_), .A3(new_n592_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  AND2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n941_), .B2(new_n942_), .ZN(G1354gat));
  AND2_X1   g744(.A1(new_n911_), .A2(new_n592_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G218gat), .B1(new_n946_), .B2(new_n482_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n658_), .A2(G218gat), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n947_), .B1(new_n946_), .B2(new_n948_), .ZN(G1355gat));
endmodule


