//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT6), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(KEYINPUT68), .A3(new_n206_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT7), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G85gat), .B(G92gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT8), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n212_), .B2(new_n207_), .ZN(new_n217_));
  OAI22_X1  g016(.A1(new_n213_), .A2(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n209_), .A2(new_n210_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(KEYINPUT64), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(G106gat), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n219_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G85gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT9), .B1(new_n229_), .B2(G92gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G85gat), .ZN(new_n233_));
  INV_X1    g032(.A(G92gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT67), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n236_));
  MUX2_X1   g035(.A(KEYINPUT67), .B(new_n235_), .S(new_n236_), .Z(new_n237_));
  OR2_X1    g036(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(new_n240_), .B2(KEYINPUT9), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n237_), .A3(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n227_), .A2(new_n228_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n228_), .B1(new_n227_), .B2(new_n242_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n218_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G57gat), .B(G64gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G78gat), .Z(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n245_), .A2(new_n252_), .ZN(new_n254_));
  OAI211_X1 g053(.A(G230gat), .B(G233gat), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT70), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT12), .B1(new_n245_), .B2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n245_), .A2(new_n252_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n245_), .A2(KEYINPUT71), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(new_n218_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n260_), .A2(KEYINPUT12), .A3(new_n262_), .A4(new_n252_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n256_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G176gat), .B(G204gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT73), .ZN(new_n268_));
  XOR2_X1   g067(.A(G120gat), .B(G148gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n270_), .B(new_n271_), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n255_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n255_), .A2(new_n275_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n265_), .A3(new_n277_), .A4(new_n272_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT13), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n274_), .B(new_n278_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n272_), .B1(new_n256_), .B2(new_n265_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n278_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n279_), .A2(new_n280_), .ZN(new_n285_));
  OAI22_X1  g084(.A1(new_n282_), .A2(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G29gat), .B(G36gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G43gat), .B(G50gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n218_), .B(new_n290_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT75), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(KEYINPUT15), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n260_), .A2(new_n262_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G232gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT34), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT35), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n297_), .A2(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n292_), .A2(new_n303_), .A3(new_n294_), .A4(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G190gat), .B(G218gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT36), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n308_), .A2(KEYINPUT36), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n302_), .A2(new_n311_), .A3(new_n304_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT37), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT37), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G231gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n252_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G8gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(G15gat), .A2(G22gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G15gat), .A2(G22gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G1gat), .A2(G8gat), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n324_), .A2(new_n325_), .B1(KEYINPUT14), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n323_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n320_), .B(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G155gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(G183gat), .B(G211gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT17), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n334_), .A2(new_n335_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n329_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n336_), .B2(new_n329_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n339_), .B(KEYINPUT78), .Z(new_n340_));
  NOR3_X1   g139(.A1(new_n287_), .A2(new_n318_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G141gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT80), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G169gat), .B(G197gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G229gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n328_), .A2(new_n290_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT79), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n328_), .A2(new_n351_), .A3(new_n290_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n328_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n293_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n328_), .A2(new_n290_), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n347_), .B(new_n357_), .C1(new_n350_), .C2(new_n352_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n346_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n353_), .A2(new_n348_), .A3(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n350_), .A2(new_n352_), .B1(new_n293_), .B2(new_n354_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n361_), .B(new_n345_), .C1(new_n348_), .C2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n356_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n366_), .A2(KEYINPUT81), .A3(new_n361_), .A4(new_n345_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  AND2_X1   g169(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n371_));
  NOR2_X1   g170(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT87), .B(new_n370_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n375_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT1), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT85), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n383_), .A2(new_n390_), .A3(KEYINPUT1), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G141gat), .B(G148gat), .Z(new_n393_));
  AOI22_X1  g192(.A1(new_n382_), .A2(new_n386_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G204gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT89), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G204gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n400_), .A3(G197gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT91), .B1(new_n397_), .B2(G197gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT89), .B(G204gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(G197gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G211gat), .B(G218gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT21), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n404_), .A2(new_n407_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n409_), .ZN(new_n415_));
  INV_X1    g214(.A(G197gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n398_), .A2(new_n400_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n409_), .B1(G197gat), .B2(G204gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT90), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n421_), .A3(new_n418_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n412_), .B1(new_n415_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G228gat), .ZN(new_n425_));
  INV_X1    g224(.A(G233gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n396_), .A2(new_n424_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n402_), .B1(new_n405_), .B2(G197gat), .ZN(new_n430_));
  AND4_X1   g229(.A1(new_n406_), .A2(new_n398_), .A3(new_n400_), .A4(G197gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n409_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n408_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n422_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n421_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n411_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT92), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n423_), .A2(new_n432_), .A3(new_n408_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT92), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n411_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n396_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n443_));
  INV_X1    g242(.A(new_n427_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n396_), .ZN(new_n446_));
  AOI211_X1 g245(.A(KEYINPUT92), .B(new_n412_), .C1(new_n415_), .C2(new_n423_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n440_), .B1(new_n439_), .B2(new_n411_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT93), .B1(new_n449_), .B2(new_n427_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n429_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n382_), .A2(new_n386_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n392_), .A2(new_n393_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT28), .B1(new_n456_), .B2(KEYINPUT29), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT28), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n394_), .A2(new_n458_), .A3(new_n395_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT88), .ZN(new_n461_));
  XOR2_X1   g260(.A(G22gat), .B(G50gat), .Z(new_n462_));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n463_), .A3(new_n459_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n443_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n449_), .A2(KEYINPUT93), .A3(new_n427_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n452_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n470_), .A2(KEYINPUT95), .A3(new_n471_), .A4(new_n429_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n453_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n471_), .B(new_n429_), .C1(new_n445_), .C2(new_n450_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n467_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n471_), .B1(new_n470_), .B2(new_n429_), .ZN(new_n478_));
  AOI211_X1 g277(.A(new_n452_), .B(new_n428_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n473_), .A2(new_n476_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT19), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G183gat), .A2(G190gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT23), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT96), .B1(G183gat), .B2(G190gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G169gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G183gat), .A2(G190gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT23), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(new_n485_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n494_), .B2(new_n485_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT96), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n499_));
  AND2_X1   g298(.A1(G169gat), .A2(G176gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G183gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT25), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(G183gat), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G190gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT26), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT26), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G190gat), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n501_), .B1(new_n506_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G169gat), .ZN(new_n513_));
  INV_X1    g312(.A(G176gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT24), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n486_), .A2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n492_), .A2(new_n498_), .B1(new_n512_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT20), .B1(new_n424_), .B2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n503_), .A2(new_n505_), .A3(new_n508_), .A4(new_n510_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT82), .B1(new_n499_), .B2(new_n500_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT82), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G169gat), .A2(G176gat), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n515_), .A2(new_n522_), .A3(KEYINPUT24), .A4(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n521_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n520_), .A2(new_n521_), .A3(new_n524_), .A4(KEYINPUT83), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n517_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n496_), .A2(new_n491_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n437_), .A2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n484_), .B1(new_n519_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT20), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n437_), .B2(new_n531_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n484_), .B1(new_n424_), .B2(new_n518_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G8gat), .B(G36gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT18), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G64gat), .B(G92gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT32), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n533_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n484_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n438_), .A2(new_n441_), .A3(new_n518_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(new_n535_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n519_), .A2(new_n532_), .A3(new_n484_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n549_), .B2(new_n543_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G127gat), .B(G134gat), .Z(new_n551_));
  XOR2_X1   g350(.A(G113gat), .B(G120gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n456_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n394_), .A2(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G225gat), .A2(G233gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT99), .B(KEYINPUT4), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(KEYINPUT4), .A3(new_n556_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n555_), .A2(KEYINPUT98), .A3(new_n556_), .A4(KEYINPUT4), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n559_), .B1(new_n566_), .B2(new_n558_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G1gat), .B(G29gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(G85gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT0), .B(G57gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n573_), .B(new_n559_), .C1(new_n566_), .C2(new_n558_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n550_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n567_), .A2(KEYINPUT33), .A3(new_n571_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT33), .B1(new_n567_), .B2(new_n571_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n533_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT97), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n533_), .A2(new_n537_), .A3(new_n581_), .A4(new_n542_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n533_), .A2(new_n537_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n541_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n566_), .A2(new_n558_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT100), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n573_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n586_), .B2(KEYINPUT100), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n585_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n575_), .B1(new_n578_), .B2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT94), .B(new_n477_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n482_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n579_), .A2(KEYINPUT27), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n541_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT101), .B(new_n541_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n542_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(KEYINPUT97), .B2(new_n579_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n604_), .B2(new_n582_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n572_), .A2(new_n574_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n476_), .A2(new_n453_), .A3(new_n467_), .A4(new_n472_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n467_), .B1(new_n453_), .B2(new_n474_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(KEYINPUT94), .ZN(new_n612_));
  INV_X1    g411(.A(new_n593_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G71gat), .B(G99gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(G43gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G227gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n616_), .B(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n531_), .B(KEYINPUT30), .Z(new_n621_));
  INV_X1    g420(.A(KEYINPUT84), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n620_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n553_), .B(KEYINPUT31), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n625_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n594_), .A2(new_n614_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n607_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n600_), .A2(new_n605_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n482_), .A2(new_n635_), .A3(new_n593_), .A4(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n369_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n341_), .A2(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n639_), .A2(G1gat), .A3(new_n608_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT38), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n480_), .A2(new_n481_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n593_), .A3(new_n610_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n572_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n567_), .A2(KEYINPUT33), .A3(new_n571_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n589_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n558_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n649_), .B(new_n561_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n582_), .B(new_n604_), .C1(new_n652_), .C2(new_n587_), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n647_), .A2(new_n653_), .B1(new_n608_), .B2(new_n550_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n633_), .B1(new_n643_), .B2(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n600_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n482_), .B2(new_n593_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n637_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT103), .A3(new_n313_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT103), .B1(new_n658_), .B2(new_n313_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n287_), .A2(new_n340_), .A3(new_n369_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n607_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G1gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n641_), .A2(new_n664_), .ZN(G1324gat));
  XNOR2_X1  g464(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n666_));
  INV_X1    g465(.A(new_n636_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n662_), .B(new_n667_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G8gat), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT39), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT39), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n639_), .A2(G8gat), .A3(new_n636_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n666_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n673_), .B(new_n666_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1325gat));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n632_), .A3(new_n662_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n632_), .A2(new_n618_), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n679_), .A2(new_n680_), .B1(new_n639_), .B2(new_n681_), .ZN(G1326gat));
  INV_X1    g481(.A(new_n643_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n639_), .A2(G22gat), .A3(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n661_), .A2(new_n643_), .A3(new_n662_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(G22gat), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n313_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n340_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n287_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n638_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n607_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n340_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n287_), .A2(new_n696_), .A3(new_n369_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT43), .B(new_n317_), .C1(new_n634_), .C2(new_n637_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n658_), .B2(new_n318_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n697_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n607_), .A2(G29gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n695_), .B1(new_n705_), .B2(new_n706_), .ZN(G1328gat));
  NOR3_X1   g506(.A1(new_n693_), .A2(G36gat), .A3(new_n636_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT45), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n703_), .A2(new_n667_), .A3(new_n704_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n710_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT106), .B1(new_n710_), .B2(G36gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI221_X1 g514(.A(new_n709_), .B1(KEYINPUT107), .B2(KEYINPUT46), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND3_X1  g516(.A1(new_n705_), .A2(G43gat), .A3(new_n632_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n693_), .B2(new_n633_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g521(.A1(new_n693_), .A2(G50gat), .A3(new_n683_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n703_), .A2(new_n643_), .A3(new_n704_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G50gat), .B1(new_n724_), .B2(new_n725_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT109), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n723_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1331gat));
  INV_X1    g531(.A(G57gat), .ZN(new_n733_));
  AND4_X1   g532(.A1(new_n661_), .A2(new_n696_), .A3(new_n369_), .A4(new_n287_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n607_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n281_), .A2(new_n286_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n318_), .A2(new_n737_), .A3(new_n340_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n368_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(G57gat), .A3(new_n608_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n735_), .A2(new_n736_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n735_), .B2(new_n741_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1332gat));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n734_), .A2(new_n667_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G64gat), .ZN(new_n747_));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT48), .B(new_n748_), .C1(new_n734_), .C2(new_n667_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n667_), .A2(new_n748_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n747_), .A2(new_n749_), .B1(new_n740_), .B2(new_n750_), .ZN(G1333gat));
  NAND2_X1  g550(.A1(new_n734_), .A2(new_n632_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G71gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G71gat), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n633_), .A2(G71gat), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT111), .Z(new_n757_));
  OAI22_X1  g556(.A1(new_n754_), .A2(new_n755_), .B1(new_n740_), .B2(new_n757_), .ZN(G1334gat));
  OR3_X1    g557(.A1(new_n740_), .A2(G78gat), .A3(new_n683_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n734_), .A2(new_n643_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G78gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G78gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n737_), .A2(new_n691_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n739_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n233_), .B1(new_n766_), .B2(new_n608_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n737_), .A2(new_n696_), .A3(new_n368_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n658_), .A2(new_n318_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT43), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n658_), .A2(new_n699_), .A3(new_n318_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n769_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n607_), .A2(new_n229_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n767_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT112), .Z(G1336gat));
  OAI21_X1  g576(.A(G92gat), .B1(new_n774_), .B2(new_n636_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n766_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n234_), .A3(new_n667_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT113), .Z(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n774_), .B2(new_n633_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n633_), .B1(new_n225_), .B2(new_n222_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g586(.A(new_n643_), .B(new_n768_), .C1(new_n698_), .C2(new_n700_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  OAI21_X1  g588(.A(G106gat), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT114), .B1(new_n773_), .B2(new_n643_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT52), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(KEYINPUT114), .A3(new_n643_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n789_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .A4(G106gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n779_), .A2(new_n203_), .A3(new_n643_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n801_), .A3(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  AOI21_X1  g602(.A(new_n346_), .B1(new_n362_), .B2(new_n348_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n357_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n348_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(new_n359_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n278_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n264_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n265_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n259_), .A2(new_n263_), .A3(KEYINPUT55), .A4(new_n264_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n273_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n273_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n808_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT58), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n273_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n815_), .B(new_n272_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT116), .B(new_n821_), .C1(new_n824_), .C2(new_n808_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n820_), .A2(new_n318_), .A3(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n368_), .A2(new_n278_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n807_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n690_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT57), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  AOI211_X1 g633(.A(KEYINPUT115), .B(new_n690_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n826_), .B(new_n831_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n340_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n737_), .A2(new_n369_), .A3(new_n317_), .A4(new_n696_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  NOR4_X1   g641(.A1(new_n643_), .A2(new_n633_), .A3(new_n667_), .A4(new_n608_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n831_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n826_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n826_), .B(KEYINPUT117), .C1(new_n834_), .C2(new_n835_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n696_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n840_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n843_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n845_), .B(new_n368_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G113gat), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n844_), .A2(G113gat), .A3(new_n369_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1340gat));
  OAI211_X1 g657(.A(new_n845_), .B(new_n287_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(G120gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n844_), .ZN(new_n861_));
  INV_X1    g660(.A(G120gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(new_n737_), .B2(KEYINPUT60), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n861_), .B(new_n863_), .C1(KEYINPUT60), .C2(new_n862_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(G1341gat));
  OAI211_X1 g664(.A(new_n845_), .B(new_n696_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G127gat), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n844_), .A2(G127gat), .A3(new_n340_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1342gat));
  OAI211_X1 g668(.A(new_n845_), .B(new_n318_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G134gat), .ZN(new_n871_));
  OR3_X1    g670(.A1(new_n844_), .A2(G134gat), .A3(new_n313_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1343gat));
  AOI21_X1  g672(.A(new_n840_), .B1(new_n340_), .B2(new_n836_), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n683_), .A2(new_n608_), .A3(new_n667_), .A4(new_n632_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n368_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n287_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n842_), .A2(new_n875_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT118), .B1(new_n882_), .B2(new_n340_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n877_), .A2(new_n884_), .A3(new_n696_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n883_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1346gat));
  OR3_X1    g688(.A1(new_n882_), .A2(G162gat), .A3(new_n313_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G162gat), .B1(new_n882_), .B2(new_n317_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1347gat));
  NAND2_X1  g691(.A1(new_n667_), .A2(new_n635_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT119), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n643_), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n368_), .B(new_n895_), .C1(new_n851_), .C2(new_n840_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n513_), .B1(new_n897_), .B2(KEYINPUT62), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(KEYINPUT62), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n896_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT22), .B(G169gat), .Z(new_n902_));
  OAI22_X1  g701(.A1(new_n900_), .A2(new_n901_), .B1(new_n896_), .B2(new_n902_), .ZN(G1348gat));
  NAND2_X1  g702(.A1(new_n287_), .A2(G176gat), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n874_), .A2(new_n643_), .A3(new_n894_), .A4(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n895_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n852_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n287_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n908_), .B2(new_n514_), .ZN(G1349gat));
  NOR2_X1   g708(.A1(new_n894_), .A2(new_n340_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n842_), .A2(new_n683_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n842_), .A2(KEYINPUT122), .A3(new_n683_), .A4(new_n910_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n502_), .A3(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n340_), .A2(new_n506_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n895_), .B(new_n916_), .C1(new_n851_), .C2(new_n840_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT121), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(KEYINPUT121), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1350gat));
  NAND2_X1  g720(.A1(new_n690_), .A2(new_n511_), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT123), .Z(new_n923_));
  NAND2_X1  g722(.A1(new_n907_), .A2(new_n923_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n852_), .A2(new_n317_), .A3(new_n906_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n507_), .B2(new_n925_), .ZN(G1351gat));
  NAND3_X1  g725(.A1(new_n643_), .A2(new_n633_), .A3(new_n608_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n667_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n842_), .A2(new_n368_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(KEYINPUT125), .B1(new_n933_), .B2(new_n416_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n874_), .A2(new_n931_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n935_), .A2(new_n936_), .A3(G197gat), .A4(new_n368_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n842_), .A2(G197gat), .A3(new_n368_), .A4(new_n932_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(KEYINPUT126), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n934_), .A2(new_n937_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n933_), .A2(new_n416_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n937_), .A2(new_n939_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n940_), .A2(new_n943_), .ZN(G1352gat));
  NAND2_X1  g743(.A1(new_n935_), .A2(new_n287_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n405_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n397_), .B2(new_n945_), .ZN(G1353gat));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n948_));
  INV_X1    g747(.A(G211gat), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n935_), .B(new_n696_), .C1(new_n948_), .C2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n949_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1354gat));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953_));
  INV_X1    g752(.A(G218gat), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n935_), .A2(new_n954_), .A3(new_n690_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n954_), .B1(new_n935_), .B2(new_n318_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n953_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n957_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n959_), .A2(new_n955_), .A3(KEYINPUT127), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n960_), .ZN(G1355gat));
endmodule


