//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_, new_n982_;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(G15gat), .ZN(new_n202_));
  INV_X1    g001(.A(G22gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  INV_X1    g004(.A(G8gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n208_), .A2(new_n209_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G29gat), .B(G36gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n217_), .A2(KEYINPUT15), .A3(new_n219_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n217_), .B2(new_n219_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n221_), .B(new_n222_), .C1(new_n213_), .C2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n222_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n212_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n220_), .B1(new_n229_), .B2(new_n210_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n220_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n211_), .A2(new_n212_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G113gat), .B(G141gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT74), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G169gat), .B(G197gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n227_), .A2(new_n233_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G78gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  INV_X1    g043(.A(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G57gat), .ZN(new_n246_));
  INV_X1    g045(.A(G57gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G64gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n243_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT66), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(new_n243_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G85gat), .B(G92gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT8), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT65), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  OR3_X1    g062(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n260_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT65), .A3(new_n258_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  INV_X1    g068(.A(G85gat), .ZN(new_n270_));
  INV_X1    g069(.A(G92gat), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT9), .ZN(new_n272_));
  XOR2_X1   g071(.A(G85gat), .B(G92gat), .Z(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(KEYINPUT9), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT10), .B(G99gat), .Z(new_n276_));
  INV_X1    g075(.A(G106gat), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT10), .B(G99gat), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n279_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n269_), .B(new_n274_), .C1(new_n278_), .C2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n258_), .A2(KEYINPUT65), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n260_), .B(new_n282_), .C1(new_n263_), .C2(new_n266_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n268_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n256_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n286_));
  INV_X1    g085(.A(new_n252_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT12), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n285_), .A2(new_n286_), .B1(new_n284_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n256_), .B2(new_n284_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT67), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n253_), .A2(new_n255_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(new_n283_), .A3(new_n281_), .A4(new_n268_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n296_), .B2(new_n291_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n290_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n285_), .A2(new_n296_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n291_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT5), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G176gat), .B(G204gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n298_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n292_), .A2(KEYINPUT67), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n296_), .A2(new_n294_), .A3(new_n291_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n312_), .A2(new_n290_), .B1(new_n300_), .B2(new_n299_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT68), .A3(new_n306_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n313_), .A2(new_n306_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n315_), .A2(KEYINPUT13), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT13), .B1(new_n315_), .B2(new_n316_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G22gat), .B(G50gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT28), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT84), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT2), .ZN(new_n332_));
  AOI211_X1 g131(.A(new_n325_), .B(new_n326_), .C1(new_n330_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G155gat), .ZN(new_n334_));
  INV_X1    g133(.A(G162gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT1), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT82), .B1(new_n336_), .B2(new_n325_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n324_), .C1(new_n326_), .C2(KEYINPUT1), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n324_), .A2(KEYINPUT1), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n329_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n331_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n342_), .A2(KEYINPUT83), .A3(new_n345_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n333_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n323_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n330_), .A2(new_n332_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n326_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n324_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n324_), .B1(new_n326_), .B2(KEYINPUT1), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n340_), .B1(new_n356_), .B2(KEYINPUT82), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n347_), .B(new_n344_), .C1(new_n357_), .C2(new_n339_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT83), .B1(new_n342_), .B2(new_n345_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n355_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n360_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n322_), .B1(new_n352_), .B2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n350_), .A2(new_n323_), .A3(new_n351_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT28), .B1(new_n360_), .B2(KEYINPUT29), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n321_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G197gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(G204gat), .ZN(new_n368_));
  INV_X1    g167(.A(G204gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G197gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G218gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G211gat), .ZN(new_n379_));
  INV_X1    g178(.A(G211gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G218gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT87), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n374_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n369_), .A2(G197gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT86), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n368_), .A2(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n370_), .B(KEYINPUT85), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n373_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n375_), .A2(new_n376_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n379_), .A2(new_n381_), .A3(new_n376_), .ZN(new_n393_));
  OAI22_X1  g192(.A1(new_n392_), .A2(new_n393_), .B1(KEYINPUT21), .B2(new_n371_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n384_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n397_), .A3(new_n395_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT88), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT89), .Z(new_n405_));
  NAND4_X1  g204(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n366_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n399_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n408_), .A2(KEYINPUT90), .ZN(new_n409_));
  INV_X1    g208(.A(new_n405_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n397_), .B1(new_n400_), .B2(new_n395_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n383_), .A2(new_n377_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n367_), .A2(G204gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT85), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n370_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n386_), .A2(new_n414_), .A3(new_n388_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT21), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n392_), .A2(new_n393_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n412_), .A2(new_n418_), .B1(new_n419_), .B2(new_n374_), .ZN(new_n420_));
  AOI211_X1 g219(.A(new_n398_), .B(new_n420_), .C1(new_n360_), .C2(KEYINPUT29), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n410_), .B1(new_n411_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n407_), .B1(new_n409_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT92), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n411_), .B2(new_n421_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n399_), .A2(KEYINPUT91), .A3(new_n401_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n404_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n408_), .A2(new_n365_), .A3(new_n362_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n424_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n408_), .A2(new_n365_), .A3(new_n362_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n426_), .A2(new_n427_), .A3(new_n404_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT92), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n423_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(G127gat), .B(G134gat), .Z(new_n435_));
  XOR2_X1   g234(.A(G113gat), .B(G120gat), .Z(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n360_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n437_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(new_n355_), .C1(new_n359_), .C2(new_n358_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G85gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n360_), .A2(new_n449_), .A3(new_n437_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT97), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n360_), .A2(new_n452_), .A3(new_n449_), .A4(new_n437_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n438_), .A2(KEYINPUT4), .A3(new_n442_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n439_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n448_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT99), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n451_), .A2(new_n453_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(new_n439_), .A3(new_n455_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT99), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n448_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT25), .B(G183gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT26), .B(G190gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G169gat), .A2(G176gat), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n464_), .A2(new_n465_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n470_));
  INV_X1    g269(.A(G169gat), .ZN(new_n471_));
  INV_X1    g270(.A(G176gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G183gat), .A2(G190gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT93), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n478_), .A2(KEYINPUT93), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n469_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n468_), .B(KEYINPUT77), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT22), .B(G169gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n472_), .B2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n476_), .A2(new_n477_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n486_), .B1(G183gat), .B2(G190gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT94), .B1(new_n489_), .B2(new_n395_), .ZN(new_n490_));
  INV_X1    g289(.A(G190gat), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n491_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n491_), .A2(KEYINPUT76), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(KEYINPUT26), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT75), .B(G183gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n483_), .A2(new_n466_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n478_), .A2(KEYINPUT78), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n478_), .A2(KEYINPUT78), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n491_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n483_), .B1(new_n486_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(G176gat), .B1(new_n471_), .B2(KEYINPUT22), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT22), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT79), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT79), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT22), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n471_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n506_), .B1(new_n511_), .B2(KEYINPUT80), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(KEYINPUT80), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n505_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n503_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n395_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n486_), .A2(new_n517_), .A3(new_n473_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n479_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n519_), .A2(new_n469_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n420_), .A3(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n490_), .A2(new_n516_), .A3(KEYINPUT20), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G226gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT19), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n489_), .A2(new_n395_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n420_), .A2(new_n503_), .A3(new_n514_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT20), .A4(new_n525_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT96), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G8gat), .B(G36gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n527_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n459_), .A2(new_n440_), .A3(new_n455_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n447_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n438_), .A2(KEYINPUT98), .A3(new_n439_), .A4(new_n442_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n540_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT33), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n540_), .A2(new_n546_), .A3(KEYINPUT33), .A4(new_n541_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n463_), .A2(new_n539_), .A3(new_n549_), .A4(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT100), .B1(new_n527_), .B2(new_n530_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n553_), .B(KEYINPUT20), .C1(new_n489_), .C2(new_n395_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n516_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n520_), .A2(new_n420_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(KEYINPUT20), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n525_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT20), .A4(new_n526_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT32), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n536_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT100), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n552_), .A2(new_n562_), .B1(new_n564_), .B2(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n547_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n541_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n434_), .A2(new_n551_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n515_), .B(KEYINPUT30), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT81), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G71gat), .B(G99gat), .ZN(new_n572_));
  INV_X1    g371(.A(G43gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G227gat), .A2(G233gat), .ZN(new_n575_));
  INV_X1    g374(.A(G15gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n574_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n570_), .B(KEYINPUT81), .Z(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n578_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n437_), .B(KEYINPUT31), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT27), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n538_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n558_), .A2(new_n559_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n536_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n584_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT102), .B1(new_n566_), .B2(new_n567_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n540_), .A2(new_n546_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n447_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n547_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n590_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n569_), .B(new_n583_), .C1(new_n434_), .C2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n582_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n581_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n590_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n591_), .A2(new_n595_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n599_), .A2(new_n434_), .A3(new_n600_), .A4(new_n601_), .ZN(new_n602_));
  AOI211_X1 g401(.A(new_n240_), .B(new_n320_), .C1(new_n597_), .C2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT35), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n268_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n225_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n284_), .A2(new_n220_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT70), .B(new_n607_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n231_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n226_), .A2(new_n284_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(KEYINPUT35), .A4(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n613_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT70), .B1(new_n616_), .B2(new_n607_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT71), .ZN(new_n619_));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT69), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT36), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n623_), .B(KEYINPUT36), .Z(new_n626_));
  OAI21_X1  g425(.A(new_n626_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT70), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(new_n624_), .A3(new_n614_), .A4(new_n611_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(KEYINPUT37), .B(new_n625_), .C1(new_n632_), .C2(new_n619_), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT72), .B(KEYINPUT37), .Z(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n213_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n252_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n287_), .ZN(new_n642_));
  XOR2_X1   g441(.A(G127gat), .B(G155gat), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT16), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT17), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(new_n642_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n640_), .A2(new_n256_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n639_), .A2(new_n295_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n646_), .B(KEYINPUT17), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n637_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n603_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n601_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n205_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n632_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n597_), .B2(new_n602_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n320_), .A2(new_n654_), .A3(new_n240_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n205_), .B1(new_n664_), .B2(new_n657_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n660_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n659_), .B2(new_n658_), .ZN(G1324gat));
  NAND3_X1  g466(.A1(new_n656_), .A2(new_n206_), .A3(new_n590_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n590_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(G8gat), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT39), .B(new_n206_), .C1(new_n664_), .C2(new_n590_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1325gat));
  AOI21_X1  g474(.A(new_n576_), .B1(new_n664_), .B2(new_n599_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT41), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n656_), .A2(new_n576_), .A3(new_n599_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1326gat));
  NOR3_X1   g478(.A1(new_n428_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT92), .B1(new_n431_), .B2(new_n432_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n409_), .A2(new_n422_), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n680_), .A2(new_n681_), .B1(new_n682_), .B2(new_n407_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n203_), .B1(new_n664_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n656_), .A2(new_n203_), .A3(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(new_n654_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n632_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n603_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n657_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n320_), .A2(new_n689_), .A3(new_n240_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT43), .B(new_n636_), .C1(new_n597_), .C2(new_n602_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n460_), .A2(new_n461_), .A3(new_n448_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n461_), .B1(new_n460_), .B2(new_n448_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n539_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n549_), .A2(new_n550_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n568_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n583_), .B1(new_n700_), .B2(new_n683_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n434_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n602_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n695_), .B1(new_n703_), .B2(new_n637_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n693_), .B1(new_n694_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n693_), .C1(new_n694_), .C2(new_n704_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n657_), .A2(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n692_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n590_), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n600_), .A2(G36gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n691_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT45), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n691_), .A2(new_n717_), .A3(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n713_), .A2(new_n719_), .A3(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  NAND4_X1  g523(.A1(new_n707_), .A2(G43gat), .A3(new_n599_), .A4(new_n708_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n691_), .A2(new_n599_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n573_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g528(.A(G50gat), .B1(new_n691_), .B2(new_n683_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n683_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n709_), .B2(new_n731_), .ZN(G1331gat));
  NAND2_X1  g531(.A1(new_n703_), .A2(new_n240_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(KEYINPUT104), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n319_), .B1(new_n733_), .B2(KEYINPUT104), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n655_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n247_), .A3(new_n657_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n240_), .A2(new_n649_), .A3(new_n653_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n319_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n662_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT105), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n662_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n742_), .A2(new_n657_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n738_), .B1(new_n247_), .B2(new_n745_), .ZN(G1332gat));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n245_), .A3(new_n590_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n590_), .A3(new_n744_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(G64gat), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n748_), .B2(G64gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n737_), .A2(new_n753_), .A3(new_n599_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n742_), .A2(new_n599_), .A3(new_n744_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G71gat), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n755_), .A3(G71gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1334gat));
  NOR2_X1   g558(.A1(new_n434_), .A2(G78gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n736_), .A2(new_n655_), .A3(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n742_), .A2(new_n683_), .A3(new_n744_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G78gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT107), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1335gat));
  NAND3_X1  g569(.A1(new_n734_), .A2(new_n690_), .A3(new_n735_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n657_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n320_), .A2(new_n654_), .A3(new_n240_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n694_), .B2(new_n704_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT108), .Z(new_n777_));
  NOR2_X1   g576(.A1(new_n601_), .A2(new_n270_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT109), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n773_), .B1(new_n777_), .B2(new_n779_), .ZN(G1336gat));
  AOI21_X1  g579(.A(G92gat), .B1(new_n772_), .B2(new_n590_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n600_), .A2(new_n271_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n777_), .B2(new_n782_), .ZN(G1337gat));
  NAND2_X1  g582(.A1(new_n599_), .A2(new_n276_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n771_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n787_));
  OAI21_X1  g586(.A(G99gat), .B1(new_n776_), .B2(new_n583_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT51), .A4(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n787_), .A2(KEYINPUT51), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(KEYINPUT51), .ZN(new_n791_));
  INV_X1    g590(.A(new_n788_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n790_), .B(new_n791_), .C1(new_n792_), .C2(new_n785_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n789_), .A2(new_n793_), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n772_), .A2(new_n277_), .A3(new_n683_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n683_), .B(new_n775_), .C1(new_n694_), .C2(new_n704_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G106gat), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n796_), .A3(G106gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n795_), .B(new_n801_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1339gat));
  AOI21_X1  g604(.A(new_n739_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n315_), .A2(new_n316_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT13), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n315_), .A2(KEYINPUT13), .A3(new_n316_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n806_), .A2(new_n809_), .A3(new_n810_), .A4(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT113), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n319_), .A2(new_n810_), .A3(new_n814_), .A4(new_n806_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n806_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT112), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n813_), .A2(new_n815_), .A3(new_n818_), .A4(new_n819_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n298_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n286_), .B1(new_n608_), .B2(new_n295_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n289_), .A2(new_n284_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n296_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT114), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n826_), .A2(new_n830_), .A3(new_n296_), .A4(new_n827_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n300_), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n312_), .A2(KEYINPUT55), .A3(new_n290_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n825_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n305_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT115), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n834_), .A2(new_n837_), .A3(KEYINPUT56), .A4(new_n305_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n834_), .A2(new_n305_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n836_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n221_), .B(new_n228_), .C1(new_n213_), .C2(new_n226_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n237_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n222_), .B1(new_n232_), .B2(new_n230_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n227_), .A2(new_n233_), .A3(new_n237_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n842_), .A2(KEYINPUT58), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n637_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n842_), .B2(new_n849_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT117), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n240_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n305_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n305_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n848_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n807_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n862_), .B2(new_n632_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  AOI211_X1 g663(.A(new_n864_), .B(new_n661_), .C1(new_n859_), .C2(new_n861_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n842_), .A2(new_n849_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n852_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n637_), .A4(new_n850_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n855_), .A2(new_n866_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n823_), .B1(new_n654_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n657_), .A2(new_n599_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n434_), .A2(new_n600_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n821_), .A2(new_n822_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n868_), .A2(new_n637_), .A3(new_n850_), .ZN(new_n879_));
  AOI211_X1 g678(.A(KEYINPUT119), .B(new_n689_), .C1(new_n866_), .C2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881_));
  INV_X1    g680(.A(new_n239_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n847_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT68), .B1(new_n313_), .B2(new_n306_), .ZN(new_n884_));
  AND4_X1   g683(.A1(KEYINPUT68), .A2(new_n298_), .A3(new_n301_), .A4(new_n306_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n841_), .B2(new_n835_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n848_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n632_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n864_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n890_), .B(new_n891_), .C1(new_n851_), .C2(new_n854_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n881_), .B1(new_n892_), .B2(new_n654_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n878_), .B1(new_n880_), .B2(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n876_), .A2(KEYINPUT118), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n876_), .A2(KEYINPUT118), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n895_), .A2(new_n896_), .A3(KEYINPUT59), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n877_), .A2(new_n898_), .A3(new_n883_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G113gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n871_), .A2(new_n654_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n878_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n875_), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n903_), .A2(G113gat), .A3(new_n240_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n904_), .ZN(G1340gat));
  INV_X1    g704(.A(new_n903_), .ZN(new_n906_));
  INV_X1    g705(.A(G120gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n319_), .B2(KEYINPUT60), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n906_), .B(new_n908_), .C1(KEYINPUT60), .C2(new_n907_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n877_), .A2(new_n898_), .A3(new_n320_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n907_), .ZN(G1341gat));
  NAND3_X1  g710(.A1(new_n877_), .A2(new_n898_), .A3(new_n689_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G127gat), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n903_), .A2(G127gat), .A3(new_n654_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1342gat));
  NAND3_X1  g714(.A1(new_n877_), .A2(new_n898_), .A3(new_n637_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G134gat), .ZN(new_n917_));
  OR3_X1    g716(.A1(new_n903_), .A2(G134gat), .A3(new_n632_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1343gat));
  NOR2_X1   g718(.A1(new_n599_), .A2(new_n434_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n600_), .A3(new_n657_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n901_), .B2(new_n878_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n883_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT120), .B(G141gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1344gat));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n320_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g726(.A1(new_n922_), .A2(new_n689_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT61), .B(G155gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1346gat));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n632_), .A2(G162gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n922_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n335_), .B1(new_n922_), .B2(new_n637_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n931_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n872_), .A2(new_n636_), .A3(new_n921_), .ZN(new_n937_));
  OAI211_X1 g736(.A(KEYINPUT121), .B(new_n933_), .C1(new_n937_), .C2(new_n335_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n657_), .A2(new_n583_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n590_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n683_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n894_), .A2(new_n883_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(G169gat), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n945_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n943_), .A2(G169gat), .A3(new_n947_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n894_), .A2(new_n942_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n949_), .A2(new_n883_), .A3(new_n484_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n946_), .A2(new_n948_), .A3(new_n950_), .ZN(G1348gat));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n320_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n872_), .A2(new_n683_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n941_), .A2(new_n472_), .A3(new_n319_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n952_), .A2(new_n472_), .B1(new_n953_), .B2(new_n954_), .ZN(G1349gat));
  NAND4_X1  g754(.A1(new_n953_), .A2(new_n689_), .A3(new_n590_), .A4(new_n940_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n654_), .A2(new_n464_), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n956_), .A2(new_n495_), .B1(new_n949_), .B2(new_n957_), .ZN(G1350gat));
  NAND2_X1  g757(.A1(new_n661_), .A2(new_n465_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(KEYINPUT123), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n949_), .A2(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n894_), .A2(new_n637_), .A3(new_n942_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(G190gat), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(G1351gat));
  NAND3_X1  g763(.A1(new_n920_), .A2(new_n590_), .A3(new_n601_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n872_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n883_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g767(.A1(new_n872_), .A2(new_n319_), .A3(new_n965_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(KEYINPUT124), .B(G204gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n969_), .B(new_n970_), .ZN(G1353gat));
  AOI21_X1  g770(.A(new_n654_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n973_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n974_));
  OR3_X1    g773(.A1(new_n973_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975_));
  AOI22_X1  g774(.A1(new_n966_), .A2(new_n972_), .B1(new_n974_), .B2(new_n975_), .ZN(new_n976_));
  AND2_X1   g775(.A1(new_n966_), .A2(new_n972_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n975_), .ZN(G1354gat));
  NAND2_X1  g777(.A1(new_n966_), .A2(new_n661_), .ZN(new_n979_));
  XOR2_X1   g778(.A(KEYINPUT126), .B(G218gat), .Z(new_n980_));
  OR2_X1    g779(.A1(new_n636_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n981_), .ZN(new_n982_));
  AOI22_X1  g781(.A1(new_n979_), .A2(new_n980_), .B1(new_n966_), .B2(new_n982_), .ZN(G1355gat));
endmodule


