//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT13), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(KEYINPUT13), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT9), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n212_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT64), .B1(new_n214_), .B2(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n216_), .A2(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n208_), .A4(new_n213_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n229_), .B1(new_n230_), .B2(KEYINPUT65), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n232_), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT66), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(KEYINPUT65), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n232_), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .A4(new_n229_), .ZN(new_n238_));
  OR2_X1    g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n216_), .A2(new_n218_), .B1(new_n239_), .B2(KEYINPUT7), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n211_), .A2(new_n212_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n228_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n228_), .B(KEYINPUT67), .C1(new_n244_), .C2(new_n245_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n251_));
  XOR2_X1   g050(.A(G71gat), .B(G78gat), .Z(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n252_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT68), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n248_), .A2(new_n249_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT69), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n241_), .A2(new_n243_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT8), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n228_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n256_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT12), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n257_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n265_), .A2(new_n266_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n274_), .B2(new_n228_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n249_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n260_), .A2(new_n261_), .A3(new_n272_), .A4(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT71), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n258_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n261_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n248_), .A2(new_n249_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n283_), .B2(new_n273_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n284_), .A2(new_n260_), .A3(new_n285_), .A4(new_n272_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n279_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G120gat), .B(G148gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT5), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G176gat), .B(G204gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  NOR2_X1   g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n291_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT72), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n292_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n203_), .B(new_n204_), .C1(new_n295_), .C2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n296_), .B2(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(KEYINPUT72), .A3(new_n294_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n202_), .A4(KEYINPUT13), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G15gat), .B(G22gat), .Z(new_n304_));
  NAND2_X1  g103(.A1(G1gat), .A2(G8gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(KEYINPUT14), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT78), .ZN(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G8gat), .Z(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n311_), .A2(new_n312_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n257_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n315_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n273_), .A3(new_n313_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G183gat), .B(G211gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n322_), .A2(KEYINPUT17), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(KEYINPUT17), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n316_), .A2(new_n318_), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n256_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n269_), .A3(new_n313_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n323_), .B(KEYINPUT79), .Z(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n326_), .A2(new_n330_), .A3(KEYINPUT80), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G232gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(KEYINPUT35), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G29gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G43gat), .B(G50gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n283_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(KEYINPUT15), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n268_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(KEYINPUT35), .A3(new_n339_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n339_), .A2(KEYINPUT35), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n349_), .A3(new_n346_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G190gat), .B(G218gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT75), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G134gat), .B(G162gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT36), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT37), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT36), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n348_), .A2(new_n359_), .A3(new_n355_), .A4(new_n350_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT77), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(KEYINPUT76), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n357_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n360_), .A2(KEYINPUT76), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT37), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n303_), .A2(new_n335_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT83), .B(G190gat), .ZN(new_n370_));
  INV_X1    g169(.A(G183gat), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n370_), .A2(KEYINPUT26), .B1(KEYINPUT25), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(KEYINPUT82), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(KEYINPUT82), .B2(new_n375_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT85), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(G176gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT24), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n382_), .B1(new_n385_), .B2(new_n380_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n391_), .A2(KEYINPUT87), .B1(KEYINPUT23), .B2(new_n387_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n393_), .A3(new_n390_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n386_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G197gat), .B(G204gat), .Z(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT21), .ZN(new_n398_));
  XOR2_X1   g197(.A(G211gat), .B(G218gat), .Z(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n401_));
  INV_X1    g200(.A(G197gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(G204gat), .ZN(new_n403_));
  OAI211_X1 g202(.A(KEYINPUT21), .B(new_n403_), .C1(new_n397_), .C2(new_n401_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n397_), .A2(new_n399_), .A3(KEYINPUT21), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n387_), .A2(new_n390_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n370_), .A2(new_n371_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(KEYINPUT88), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(new_n383_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n412_), .B2(KEYINPUT88), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n396_), .A2(new_n408_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n391_), .A2(KEYINPUT87), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n387_), .A2(KEYINPUT23), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n394_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G190gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n371_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n415_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n409_), .A2(new_n410_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n380_), .B1(new_n385_), .B2(KEYINPUT99), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(KEYINPUT99), .B2(new_n385_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT25), .B(G183gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT26), .B(G190gat), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n428_), .A2(new_n429_), .B1(new_n381_), .B2(new_n380_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n407_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n418_), .A2(KEYINPUT20), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n396_), .A2(new_n417_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n407_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n424_), .A2(new_n432_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n436_), .B1(new_n440_), .B2(new_n408_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT20), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT18), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT101), .B1(new_n424_), .B2(new_n432_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n392_), .A2(new_n394_), .B1(new_n371_), .B2(new_n422_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n449_), .B(new_n431_), .C1(new_n450_), .C2(new_n415_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n448_), .A2(new_n408_), .A3(new_n451_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n379_), .A2(new_n395_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT20), .B1(new_n453_), .B2(new_n408_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n436_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n453_), .B2(new_n408_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n436_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n433_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT27), .B(new_n447_), .C1(new_n460_), .C2(new_n446_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n446_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n458_), .B1(new_n457_), .B2(new_n433_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n431_), .B1(new_n450_), .B2(new_n415_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n458_), .B1(new_n464_), .B2(new_n407_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n454_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n447_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT27), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n461_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G113gat), .B(G120gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT90), .ZN(new_n474_));
  XOR2_X1   g273(.A(G127gat), .B(G134gat), .Z(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n474_), .A2(new_n475_), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT91), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT31), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT89), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n485_), .B(G15gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT30), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n484_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(G43gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n453_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n492_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G29gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G85gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT0), .B(G57gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  NOR2_X1   g298(.A1(G155gat), .A2(G162gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT1), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G155gat), .A2(G162gat), .ZN(new_n502_));
  MUX2_X1   g301(.A(KEYINPUT1), .B(new_n501_), .S(new_n502_), .Z(new_n503_));
  NAND2_X1  g302(.A1(G141gat), .A2(G148gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT92), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G141gat), .A2(G148gat), .ZN(new_n507_));
  MUX2_X1   g306(.A(new_n506_), .B(new_n505_), .S(new_n507_), .Z(new_n508_));
  NOR2_X1   g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n502_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(new_n500_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n507_), .B(KEYINPUT3), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT2), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n517_), .A2(KEYINPUT93), .B1(G141gat), .B2(G148gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(KEYINPUT93), .B2(new_n517_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT95), .A4(new_n519_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n512_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n478_), .B(new_n481_), .C1(new_n509_), .C2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n474_), .B(new_n475_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n509_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n522_), .A2(new_n523_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n526_), .B(new_n527_), .C1(new_n528_), .C2(new_n512_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(KEYINPUT4), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT100), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n525_), .A2(KEYINPUT100), .A3(new_n529_), .A4(KEYINPUT4), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G225gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n525_), .B2(KEYINPUT4), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n525_), .A2(new_n529_), .A3(new_n535_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n499_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n540_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n499_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G228gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT96), .Z(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT29), .B1(new_n524_), .B2(new_n509_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n407_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G78gat), .B(G106gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n407_), .A3(new_n548_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT98), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n557_), .B2(new_n550_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n524_), .A2(KEYINPUT29), .A3(new_n509_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G22gat), .B(G50gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT28), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n559_), .B(new_n561_), .ZN(new_n562_));
  AND4_X1   g361(.A1(new_n555_), .A2(new_n556_), .A3(new_n558_), .A4(new_n562_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n556_), .A2(new_n562_), .B1(new_n558_), .B2(new_n555_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n472_), .A2(new_n495_), .A3(new_n546_), .A4(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n544_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n539_), .A2(new_n540_), .A3(new_n499_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n567_), .B(new_n568_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n471_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n446_), .A2(KEYINPUT32), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n455_), .B2(new_n459_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n437_), .A2(new_n442_), .A3(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT102), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n574_), .B(KEYINPUT102), .C1(new_n541_), .C2(new_n545_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n568_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n525_), .A2(new_n529_), .A3(new_n536_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n544_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n525_), .A2(KEYINPUT4), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n536_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n534_), .B2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n468_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n545_), .A2(KEYINPUT33), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n577_), .A2(new_n578_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n570_), .B1(new_n589_), .B2(new_n565_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n566_), .B1(new_n590_), .B2(new_n495_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n311_), .A2(new_n345_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT81), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n309_), .A2(new_n343_), .A3(new_n310_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G229gat), .A2(G233gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n311_), .B(new_n343_), .Z(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  AND3_X1   g401(.A1(new_n596_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n591_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n369_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n546_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(KEYINPUT103), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(KEYINPUT103), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n608_), .A2(G1gat), .A3(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT38), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n357_), .A2(new_n360_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n591_), .A2(KEYINPUT104), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT104), .B1(new_n591_), .B2(new_n616_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n303_), .A2(new_n331_), .A3(new_n605_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n609_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G1gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(new_n622_), .ZN(G1324gat));
  XNOR2_X1  g422(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n471_), .B(new_n620_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626_));
  AND4_X1   g425(.A1(KEYINPUT105), .A2(new_n625_), .A3(new_n626_), .A4(G8gat), .ZN(new_n627_));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(KEYINPUT39), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n625_), .A2(new_n630_), .B1(KEYINPUT105), .B2(new_n626_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n608_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n628_), .A3(new_n471_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n624_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n634_), .B(new_n624_), .C1(new_n627_), .C2(new_n631_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1325gat));
  NAND3_X1  g437(.A1(new_n619_), .A2(new_n495_), .A3(new_n620_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G15gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT41), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n642_), .A3(G15gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT107), .ZN(new_n644_));
  INV_X1    g443(.A(new_n495_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n633_), .B2(new_n646_), .ZN(new_n647_));
  NOR4_X1   g446(.A1(new_n608_), .A2(KEYINPUT107), .A3(G15gat), .A4(new_n645_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n641_), .A2(new_n643_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT108), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n641_), .A2(new_n652_), .A3(new_n643_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1326gat));
  OR3_X1    g453(.A1(new_n608_), .A2(G22gat), .A3(new_n565_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n565_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n619_), .A2(new_n656_), .A3(new_n620_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G22gat), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(KEYINPUT42), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(KEYINPUT42), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n659_), .B2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n335_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n303_), .A2(new_n605_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(KEYINPUT109), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n591_), .A2(new_n368_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(KEYINPUT109), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n591_), .A2(new_n368_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n663_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT44), .B(new_n663_), .C1(new_n667_), .C2(new_n669_), .ZN(new_n673_));
  AND4_X1   g472(.A1(G29gat), .A2(new_n672_), .A3(new_n612_), .A4(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n303_), .A2(new_n616_), .A3(new_n662_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n607_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n609_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n674_), .A2(new_n678_), .ZN(G1328gat));
  AOI21_X1  g478(.A(KEYINPUT110), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n471_), .A3(new_n673_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n472_), .A2(G36gat), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n677_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT45), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n677_), .A2(new_n686_), .A3(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n680_), .B1(new_n682_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n682_), .A2(new_n690_), .A3(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT111), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(G1329gat));
  NAND4_X1  g493(.A1(new_n672_), .A2(G43gat), .A3(new_n495_), .A4(new_n673_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n676_), .A2(new_n645_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(G43gat), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g497(.A1(G50gat), .A2(new_n672_), .A3(new_n656_), .A4(new_n673_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G50gat), .B1(new_n677_), .B2(new_n656_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1331gat));
  AND2_X1   g500(.A1(new_n591_), .A2(new_n605_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n702_), .A2(new_n303_), .A3(new_n662_), .A4(new_n367_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT112), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n612_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n303_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n596_), .A2(new_n599_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n602_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n596_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n710_), .A2(new_n333_), .A3(new_n711_), .A4(new_n334_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n619_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n546_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n706_), .A2(new_n715_), .ZN(G1332gat));
  INV_X1    g515(.A(G64gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n704_), .A2(new_n717_), .A3(new_n471_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719_));
  INV_X1    g518(.A(new_n714_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n471_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n721_), .B2(G64gat), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT48), .B(new_n717_), .C1(new_n720_), .C2(new_n471_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(G1333gat));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n704_), .A2(new_n725_), .A3(new_n495_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT49), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n720_), .A2(new_n495_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G71gat), .ZN(new_n729_));
  AOI211_X1 g528(.A(KEYINPUT49), .B(new_n725_), .C1(new_n720_), .C2(new_n495_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1334gat));
  NOR2_X1   g530(.A1(new_n565_), .A2(G78gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT115), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n704_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n619_), .A2(new_n656_), .A3(new_n713_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G78gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n738_), .A3(G78gat), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n737_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n734_), .B1(new_n741_), .B2(new_n742_), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n591_), .A2(new_n605_), .ZN(new_n744_));
  NOR4_X1   g543(.A1(new_n744_), .A2(new_n707_), .A3(new_n616_), .A4(new_n662_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n612_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n606_), .A2(new_n662_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n303_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n303_), .B2(new_n748_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n667_), .A2(new_n669_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n609_), .A2(G85gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT117), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n746_), .A2(G85gat), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT118), .ZN(G1336gat));
  OAI21_X1  g554(.A(G92gat), .B1(new_n751_), .B2(new_n472_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n745_), .A2(new_n210_), .A3(new_n471_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1337gat));
  NAND4_X1  g557(.A1(new_n745_), .A2(new_n495_), .A3(new_n205_), .A4(new_n207_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G99gat), .B1(new_n751_), .B2(new_n645_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT119), .B(G99gat), .C1(new_n751_), .C2(new_n645_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n745_), .A2(new_n206_), .A3(new_n656_), .ZN(new_n769_));
  OAI221_X1 g568(.A(new_n656_), .B1(new_n749_), .B2(new_n750_), .C1(new_n669_), .C2(new_n667_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G106gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g574(.A1(new_n645_), .A2(new_n656_), .A3(new_n471_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n612_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  INV_X1    g578(.A(new_n291_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n260_), .A2(new_n277_), .A3(new_n272_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n281_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n278_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n279_), .A2(new_n783_), .A3(new_n286_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT122), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n279_), .A2(KEYINPUT122), .A3(new_n783_), .A4(new_n286_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n779_), .B(new_n780_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n784_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n291_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n789_), .A2(new_n793_), .A3(KEYINPUT123), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n291_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT123), .A3(new_n779_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n593_), .A2(new_n594_), .A3(new_n598_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n602_), .B1(new_n597_), .B2(new_n595_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n711_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(new_n292_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n796_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n778_), .B1(new_n794_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n793_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n291_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n801_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n793_), .B2(KEYINPUT123), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n803_), .A2(new_n368_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT124), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n803_), .A2(new_n810_), .A3(new_n813_), .A4(new_n368_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n605_), .A2(new_n292_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n789_), .B2(new_n793_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n800_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT57), .B1(new_n819_), .B2(new_n616_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  INV_X1    g620(.A(new_n616_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n821_), .B(new_n822_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n812_), .A2(new_n814_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n331_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n712_), .B(KEYINPUT121), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n367_), .A2(new_n299_), .A3(new_n827_), .A4(new_n302_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n777_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n606_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n823_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n819_), .A2(new_n616_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n821_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n811_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n830_), .B1(new_n839_), .B2(new_n335_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n777_), .A2(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n605_), .A2(new_n834_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT125), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n843_), .B(new_n845_), .C1(new_n832_), .C2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n835_), .A2(new_n847_), .ZN(G1340gat));
  OAI211_X1 g647(.A(new_n303_), .B(new_n843_), .C1(new_n832_), .C2(new_n846_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n832_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n832_), .A2(new_n662_), .ZN(new_n855_));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n331_), .A2(new_n856_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n843_), .B(new_n858_), .C1(new_n832_), .C2(new_n846_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1342gat));
  NAND2_X1  g659(.A1(new_n832_), .A2(new_n822_), .ZN(new_n861_));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT126), .B(G134gat), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n367_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n843_), .B(new_n865_), .C1(new_n832_), .C2(new_n846_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n863_), .A2(new_n866_), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n826_), .A2(new_n831_), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n613_), .A2(new_n565_), .A3(new_n471_), .A4(new_n495_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n606_), .A3(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g670(.A1(new_n868_), .A2(new_n303_), .A3(new_n869_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g672(.A1(new_n868_), .A2(new_n662_), .A3(new_n869_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  AND2_X1   g675(.A1(new_n868_), .A2(new_n869_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n822_), .ZN(new_n878_));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n367_), .A2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT127), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n878_), .A2(new_n879_), .B1(new_n877_), .B2(new_n881_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n645_), .A2(new_n472_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n613_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n565_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n662_), .B1(new_n824_), .B2(new_n811_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n606_), .B(new_n887_), .C1(new_n888_), .C2(new_n830_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT62), .B(new_n383_), .C1(new_n889_), .C2(KEYINPUT22), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  INV_X1    g690(.A(new_n889_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT22), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G169gat), .B1(new_n889_), .B2(KEYINPUT62), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n890_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(G1348gat));
  NOR2_X1   g696(.A1(new_n840_), .A2(new_n886_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G176gat), .B1(new_n898_), .B2(new_n303_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n656_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n707_), .A2(new_n384_), .A3(new_n884_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  INV_X1    g701(.A(new_n898_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n903_), .A2(new_n428_), .A3(new_n331_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n662_), .A3(new_n885_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n371_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n903_), .B2(new_n367_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n898_), .A2(new_n429_), .A3(new_n822_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n472_), .A2(new_n495_), .A3(new_n569_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n606_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n303_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g715(.A(new_n331_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n912_), .B(new_n917_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n912_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n331_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n922_), .B2(new_n918_), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n921_), .B2(new_n367_), .ZN(new_n924_));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n912_), .A2(new_n925_), .A3(new_n822_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1355gat));
endmodule


