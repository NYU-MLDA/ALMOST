//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT78), .ZN(new_n207_));
  OR2_X1    g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(KEYINPUT1), .B2(new_n205_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n203_), .B(new_n204_), .C1(new_n207_), .C2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n203_), .A2(KEYINPUT3), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n203_), .A2(KEYINPUT3), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(new_n204_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(KEYINPUT79), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(new_n212_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n205_), .A3(new_n208_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G22gat), .B(G50gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n222_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT80), .B(KEYINPUT28), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT83), .B(G197gat), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT84), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n232_), .A3(new_n229_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT85), .B(G204gat), .Z(new_n234_));
  OAI211_X1 g033(.A(new_n231_), .B(new_n233_), .C1(G197gat), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT21), .ZN(new_n236_));
  XOR2_X1   g035(.A(G211gat), .B(G218gat), .Z(new_n237_));
  INV_X1    g036(.A(new_n228_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n238_), .A2(G204gat), .B1(new_n234_), .B2(G197gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n239_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n234_), .A2(G197gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(new_n229_), .B2(new_n228_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT86), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n247_), .A3(new_n237_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT82), .B1(new_n219_), .B2(KEYINPUT29), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G228gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G78gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n255_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT81), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n227_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264_));
  INV_X1    g063(.A(G113gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(G120gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT89), .A3(new_n219_), .ZN(new_n268_));
  INV_X1    g067(.A(G120gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n266_), .B(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n218_), .A3(new_n210_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n263_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n268_), .A2(new_n263_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n262_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n219_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n261_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G57gat), .B(G85gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT91), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n279_), .B(new_n280_), .Z(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n281_), .B(new_n282_), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n274_), .A2(new_n276_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT23), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(G183gat), .B2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT74), .B(G176gat), .Z(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT22), .B(G169gat), .Z(new_n294_));
  OAI211_X1 g093(.A(new_n291_), .B(new_n292_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n298_), .A2(new_n290_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT30), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT75), .B(KEYINPUT76), .Z(new_n308_));
  NAND2_X1  g107(.A1(G227gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G71gat), .B(G99gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G15gat), .B(G43gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n306_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n307_), .B1(new_n306_), .B2(new_n314_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n270_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n267_), .A3(new_n315_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n304_), .A2(new_n305_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n318_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n288_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n295_), .A2(new_n302_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n242_), .A2(new_n248_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT20), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(KEYINPUT20), .B(new_n336_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n331_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n340_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n249_), .A2(new_n303_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n242_), .A2(new_n332_), .A3(new_n248_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n336_), .B1(new_n347_), .B2(KEYINPUT20), .ZN(new_n348_));
  INV_X1    g147(.A(new_n339_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n344_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n330_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n343_), .A2(KEYINPUT27), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT27), .B1(new_n343_), .B2(new_n352_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n325_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n343_), .A2(new_n352_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n343_), .A2(new_n352_), .A3(KEYINPUT27), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT95), .A3(new_n359_), .ZN(new_n360_));
  AOI211_X1 g159(.A(new_n260_), .B(new_n324_), .C1(new_n355_), .C2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n353_), .A2(new_n354_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n259_), .B1(new_n363_), .B2(new_n288_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT32), .B(new_n330_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n350_), .A2(new_n351_), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n287_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n286_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n271_), .A2(new_n275_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n261_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT93), .B1(new_n285_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n261_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT93), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n283_), .B(new_n375_), .C1(new_n261_), .C2(new_n371_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n343_), .A2(new_n352_), .A3(new_n370_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n286_), .A2(new_n369_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT92), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n259_), .B(new_n368_), .C1(new_n378_), .C2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n322_), .A2(new_n323_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n362_), .B1(new_n364_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n358_), .A2(new_n288_), .A3(new_n359_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n260_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(KEYINPUT94), .A3(new_n382_), .A4(new_n381_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n361_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G120gat), .B(G148gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(new_n229_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT5), .ZN(new_n391_));
  INV_X1    g190(.A(G176gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT7), .ZN(new_n395_));
  INV_X1    g194(.A(G99gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n254_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G99gat), .A2(G106gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n397_), .A2(new_n400_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(G85gat), .A2(G92gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G85gat), .A2(G92gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT8), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT8), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(new_n409_), .A3(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n404_), .A2(KEYINPUT9), .A3(new_n405_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n405_), .A2(KEYINPUT9), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n396_), .A2(KEYINPUT10), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n396_), .A2(KEYINPUT10), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n254_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT65), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT10), .B(G99gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(G106gat), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n411_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G78gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(G57gat), .A2(G64gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT11), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G57gat), .A2(G64gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(G57gat), .A2(G64gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G57gat), .A2(G64gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT11), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n429_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n428_), .B(KEYINPUT11), .C1(new_n435_), .C2(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT12), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n427_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT12), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n408_), .A2(new_n410_), .B1(new_n420_), .B2(new_n417_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n437_), .A2(new_n438_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G230gat), .ZN(new_n446_));
  INV_X1    g245(.A(G233gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT66), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n441_), .A2(new_n445_), .A3(new_n449_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n420_), .A2(new_n414_), .A3(new_n416_), .A4(new_n415_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n403_), .A2(new_n409_), .A3(new_n406_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n409_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n444_), .B(new_n456_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT64), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT64), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n411_), .A2(new_n461_), .A3(new_n456_), .A4(new_n444_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n444_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n467_), .A2(new_n448_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n394_), .B1(new_n455_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n454_), .A3(new_n393_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n472_), .A2(KEYINPUT13), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(KEYINPUT13), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G50gat), .ZN(new_n485_));
  INV_X1    g284(.A(G29gat), .ZN(new_n486_));
  INV_X1    g285(.A(G36gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G43gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n485_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G29gat), .B(G36gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(G43gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G50gat), .A3(new_n491_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n494_), .A2(KEYINPUT15), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT15), .B1(new_n494_), .B2(new_n497_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n484_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n482_), .A2(new_n483_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n492_), .A2(new_n485_), .A3(new_n493_), .ZN(new_n502_));
  AOI21_X1  g301(.A(G50gat), .B1(new_n496_), .B2(new_n491_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n500_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n501_), .A2(new_n504_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n484_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT73), .B(G141gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT72), .B(G113gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n511_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n476_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n484_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(new_n444_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT70), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT16), .B(G183gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G211gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G127gat), .B(G155gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT17), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT71), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n526_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n523_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n539_), .A2(KEYINPUT96), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(KEYINPUT96), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT67), .B(G134gat), .ZN(new_n542_));
  INV_X1    g341(.A(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT36), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n427_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n443_), .A2(new_n504_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(KEYINPUT35), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n548_), .A2(new_n555_), .A3(new_n556_), .A4(new_n549_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n553_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n554_), .B1(new_n553_), .B2(new_n557_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n547_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n553_), .A2(new_n563_), .A3(new_n546_), .A4(new_n557_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT69), .B(new_n547_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR4_X1   g366(.A1(new_n388_), .A2(new_n540_), .A3(new_n541_), .A4(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n202_), .B1(new_n568_), .B2(new_n287_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT97), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n553_), .A2(new_n557_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n547_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT37), .A3(new_n564_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(new_n475_), .A3(new_n538_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n388_), .A2(new_n522_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n202_), .A3(new_n287_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT38), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n570_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT98), .Z(G1324gat));
  INV_X1    g382(.A(new_n355_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n360_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n478_), .B1(new_n568_), .B2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT39), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n579_), .A2(new_n478_), .A3(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g390(.A(G15gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n382_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n568_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT41), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n579_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1326gat));
  INV_X1    g396(.A(G22gat), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n598_), .B1(new_n568_), .B2(new_n260_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT42), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n579_), .A2(new_n598_), .A3(new_n260_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT99), .Z(G1327gat));
  NAND2_X1  g402(.A1(new_n384_), .A2(new_n387_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n361_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n567_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n538_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n523_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n287_), .A2(new_n486_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT101), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n614_));
  INV_X1    g413(.A(new_n609_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n606_), .B2(new_n576_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n388_), .A2(KEYINPUT43), .A3(new_n577_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n615_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n614_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n606_), .A2(new_n616_), .A3(new_n576_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT43), .B1(new_n388_), .B2(new_n577_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n609_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n624_), .A2(KEYINPUT100), .A3(KEYINPUT44), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT44), .B(new_n615_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n626_), .A2(new_n288_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n613_), .B1(new_n629_), .B2(new_n486_), .ZN(G1328gat));
  NAND3_X1  g429(.A1(new_n610_), .A2(new_n586_), .A3(new_n487_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT45), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n586_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT100), .B1(new_n624_), .B2(KEYINPUT44), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n619_), .A2(new_n614_), .A3(new_n620_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n632_), .B(KEYINPUT46), .C1(new_n636_), .C2(new_n487_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT104), .ZN(new_n638_));
  INV_X1    g437(.A(new_n586_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n624_), .B2(KEYINPUT44), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G36gat), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(KEYINPUT46), .A4(new_n632_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n638_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n632_), .B1(new_n636_), .B2(new_n487_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT102), .B(KEYINPUT46), .Z(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT103), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(KEYINPUT103), .A3(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1329gat));
  OAI211_X1 g449(.A(new_n593_), .B(new_n627_), .C1(new_n621_), .C2(new_n625_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n382_), .A2(G43gat), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n651_), .A2(G43gat), .B1(new_n610_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g453(.A(G50gat), .B1(new_n610_), .B2(new_n260_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n626_), .A2(new_n628_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n259_), .A2(new_n485_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(G1331gat));
  NOR2_X1   g457(.A1(new_n388_), .A2(new_n521_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n608_), .A2(new_n475_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n577_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT105), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(KEYINPUT105), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n287_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n566_), .A3(new_n660_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT106), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(new_n287_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n669_), .B2(G57gat), .ZN(G1332gat));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n586_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G64gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT107), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n671_), .A2(new_n674_), .A3(G64gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(KEYINPUT48), .A3(new_n675_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n664_), .A2(G64gat), .A3(new_n639_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(G1333gat));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n668_), .B2(new_n593_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT49), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n665_), .A2(new_n682_), .A3(new_n593_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1334gat));
  NAND2_X1  g485(.A1(new_n668_), .A2(new_n260_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G78gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT50), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n259_), .A2(G78gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n664_), .B2(new_n690_), .ZN(G1335gat));
  NAND3_X1  g490(.A1(new_n608_), .A2(new_n522_), .A3(new_n476_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n607_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n287_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n622_), .A2(new_n623_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n692_), .B(KEYINPUT108), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT109), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n287_), .A2(G85gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT110), .Z(new_n700_));
  AOI21_X1  g499(.A(new_n694_), .B1(new_n698_), .B2(new_n700_), .ZN(G1336gat));
  INV_X1    g500(.A(G92gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n693_), .A2(new_n586_), .A3(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n698_), .A2(new_n586_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n702_), .ZN(G1337gat));
  OAI21_X1  g504(.A(G99gat), .B1(new_n697_), .B2(new_n382_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n693_), .B(new_n593_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g508(.A1(new_n693_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G106gat), .B1(new_n697_), .B2(new_n259_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT52), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(KEYINPUT52), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g514(.A(KEYINPUT117), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n471_), .A2(new_n521_), .ZN(new_n717_));
  AND4_X1   g516(.A1(KEYINPUT111), .A2(new_n463_), .A3(new_n445_), .A4(new_n441_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n414_), .A2(new_n415_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n719_), .A2(KEYINPUT65), .A3(new_n420_), .A4(new_n416_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n423_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n439_), .B1(new_n722_), .B2(new_n411_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT12), .B1(new_n464_), .B2(new_n465_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT111), .B1(new_n725_), .B2(new_n463_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n448_), .B1(new_n718_), .B2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT112), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n448_), .C1(new_n718_), .C2(new_n726_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT113), .B1(new_n450_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n725_), .A2(new_n733_), .A3(KEYINPUT55), .A4(new_n449_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n454_), .A2(new_n731_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n728_), .A2(new_n730_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n394_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT56), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(KEYINPUT56), .A3(new_n394_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n717_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n500_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n506_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n516_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n518_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n472_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n566_), .B1(new_n741_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n745_), .B(KEYINPUT114), .ZN(new_n754_));
  INV_X1    g553(.A(new_n471_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n747_), .A2(KEYINPUT115), .A3(new_n471_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n736_), .A2(KEYINPUT56), .A3(new_n394_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT56), .B1(new_n736_), .B2(new_n394_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n758_), .B(KEYINPUT58), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(KEYINPUT116), .A3(new_n576_), .A4(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n752_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n576_), .A3(new_n764_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n521_), .B(new_n471_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n567_), .B1(new_n769_), .B2(new_n748_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n767_), .A2(new_n768_), .B1(new_n770_), .B2(KEYINPUT57), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n538_), .B1(new_n766_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n577_), .A2(new_n538_), .A3(new_n522_), .A4(new_n475_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n716_), .B1(new_n772_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n767_), .A2(new_n768_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n770_), .A2(KEYINPUT57), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n752_), .A4(new_n765_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n608_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n773_), .B(KEYINPUT54), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(KEYINPUT117), .A3(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n776_), .A2(new_n782_), .ZN(new_n783_));
  NOR4_X1   g582(.A1(new_n586_), .A2(new_n288_), .A3(new_n260_), .A4(new_n382_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n265_), .B1(new_n785_), .B2(new_n522_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(KEYINPUT59), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT119), .B1(new_n752_), .B2(new_n767_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(KEYINPUT57), .B2(new_n770_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n752_), .A2(KEYINPUT119), .A3(new_n767_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n608_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n781_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n784_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n789_), .A2(G113gat), .A3(new_n797_), .A4(new_n521_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n787_), .A2(new_n788_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT120), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n787_), .A2(new_n801_), .A3(new_n788_), .A4(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1340gat));
  INV_X1    g602(.A(new_n785_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n269_), .B1(new_n475_), .B2(KEYINPUT60), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n804_), .B(new_n805_), .C1(KEYINPUT60), .C2(new_n269_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n789_), .A2(new_n797_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n476_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n806_), .B1(new_n808_), .B2(new_n269_), .ZN(G1341gat));
  AOI21_X1  g608(.A(G127gat), .B1(new_n804_), .B2(new_n538_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n807_), .A2(G127gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n538_), .ZN(G1342gat));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n785_), .B2(new_n566_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n814_), .A2(KEYINPUT121), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(KEYINPUT121), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n576_), .A2(G134gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT122), .Z(new_n818_));
  AOI22_X1  g617(.A1(new_n815_), .A2(new_n816_), .B1(new_n807_), .B2(new_n818_), .ZN(G1343gat));
  NOR2_X1   g618(.A1(new_n593_), .A2(new_n259_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n783_), .A2(new_n287_), .A3(new_n639_), .A4(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n522_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT123), .B(G141gat), .Z(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1344gat));
  NOR2_X1   g623(.A1(new_n821_), .A2(new_n475_), .ZN(new_n825_));
  XOR2_X1   g624(.A(new_n825_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g625(.A1(new_n821_), .A2(new_n608_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT61), .B(G155gat), .Z(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(G1346gat));
  NOR3_X1   g628(.A1(new_n821_), .A2(new_n543_), .A3(new_n577_), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n821_), .A2(new_n566_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n543_), .B2(new_n831_), .ZN(G1347gat));
  AOI21_X1  g631(.A(new_n260_), .B1(new_n794_), .B2(new_n781_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n639_), .A2(new_n324_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G169gat), .B1(new_n835_), .B2(new_n522_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n835_), .A2(new_n522_), .A3(new_n294_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n837_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(G1348gat));
  NAND3_X1  g640(.A1(new_n833_), .A2(new_n476_), .A3(new_n834_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n293_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n783_), .A2(new_n259_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n639_), .A2(new_n392_), .A3(new_n475_), .A4(new_n324_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n842_), .A2(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(G1349gat));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n538_), .A3(new_n834_), .ZN(new_n847_));
  INV_X1    g646(.A(G183gat), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n639_), .A2(new_n608_), .A3(new_n296_), .A4(new_n324_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n847_), .A2(new_n848_), .B1(new_n833_), .B2(new_n849_), .ZN(G1350gat));
  OAI21_X1  g649(.A(G190gat), .B1(new_n835_), .B2(new_n577_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n833_), .A2(new_n297_), .A3(new_n834_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n566_), .B2(new_n852_), .ZN(G1351gat));
  AND3_X1   g652(.A1(new_n586_), .A2(new_n288_), .A3(new_n820_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n776_), .A2(new_n782_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT124), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n776_), .A2(new_n782_), .A3(new_n857_), .A4(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n521_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n476_), .ZN(new_n862_));
  MUX2_X1   g661(.A(new_n234_), .B(G204gat), .S(new_n862_), .Z(G1353gat));
  AOI21_X1  g662(.A(new_n608_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n859_), .A2(new_n538_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n865_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n864_), .A2(KEYINPUT125), .A3(new_n866_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT126), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n875_), .B(new_n868_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1354gat));
  INV_X1    g676(.A(G218gat), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n878_), .B(new_n577_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n859_), .A2(new_n567_), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT127), .Z(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n881_), .B2(new_n878_), .ZN(G1355gat));
endmodule


