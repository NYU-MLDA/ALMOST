//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT82), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n210_), .A3(KEYINPUT22), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT83), .B(G176gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT23), .ZN(new_n216_));
  OR2_X1    g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n216_), .A2(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n203_), .A2(new_n220_), .A3(KEYINPUT80), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n221_), .A2(new_n223_), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n225_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n231_), .A2(new_n216_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n219_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT30), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n214_), .A2(new_n218_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n202_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G113gat), .B(G120gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(new_n240_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n202_), .B(new_n245_), .C1(new_n235_), .C2(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT31), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n234_), .A2(KEYINPUT30), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n236_), .A2(new_n237_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT84), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(G71gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G99gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G15gat), .B(G43gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n248_), .B1(new_n251_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n247_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n251_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n246_), .B(new_n243_), .C1(new_n262_), .C2(new_n258_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G197gat), .B(G204gat), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  INV_X1    g067(.A(G204gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(G197gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(KEYINPUT21), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n265_), .A2(KEYINPUT21), .A3(new_n267_), .A4(new_n270_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277_));
  INV_X1    g076(.A(G141gat), .ZN(new_n278_));
  INV_X1    g077(.A(G148gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G141gat), .A2(G148gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n280_), .A2(new_n283_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G155gat), .ZN(new_n287_));
  INV_X1    g086(.A(G162gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G155gat), .A2(G162gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n293_), .A2(KEYINPUT1), .B1(new_n278_), .B2(new_n279_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n295_), .A3(new_n290_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n296_), .A3(new_n281_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n276_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(G78gat), .B1(new_n275_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n275_), .A2(new_n298_), .A3(G78gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n272_), .A2(new_n274_), .A3(KEYINPUT86), .A4(new_n273_), .ZN(new_n302_));
  INV_X1    g101(.A(G106gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G228gat), .A2(G233gat), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n300_), .A2(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n304_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G106gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n275_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n298_), .ZN(new_n311_));
  INV_X1    g110(.A(G78gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(new_n313_), .A3(new_n299_), .A4(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n307_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G22gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G50gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n292_), .A2(new_n297_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(KEYINPUT29), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n320_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n307_), .A2(new_n315_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(KEYINPUT88), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n316_), .B(KEYINPUT89), .C1(new_n307_), .C2(new_n315_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n325_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n328_), .A2(new_n330_), .A3(new_n324_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n264_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n325_), .A3(new_n331_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n324_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n321_), .A2(KEYINPUT92), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n292_), .A2(new_n340_), .A3(new_n297_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n341_), .A3(new_n245_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n321_), .A2(new_n242_), .A3(KEYINPUT92), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n245_), .A2(new_n321_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n341_), .A2(new_n245_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n340_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n343_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT4), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT93), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n344_), .A2(new_n358_), .A3(KEYINPUT4), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n351_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n348_), .B1(new_n360_), .B2(new_n345_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362_));
  INV_X1    g161(.A(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT0), .B(G57gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT97), .B1(new_n361_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n367_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n358_), .B1(new_n344_), .B2(KEYINPUT4), .ZN(new_n370_));
  AOI211_X1 g169(.A(KEYINPUT93), .B(new_n349_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n350_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n347_), .B1(new_n372_), .B2(new_n346_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n366_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n368_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT18), .B(G64gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n225_), .B1(G169gat), .B2(G176gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n227_), .B2(new_n225_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n232_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n213_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n218_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n275_), .A3(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(KEYINPUT20), .C1(new_n236_), .C2(new_n275_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT19), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT91), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n234_), .A2(new_n310_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT91), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT20), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n232_), .A2(new_n384_), .B1(new_n218_), .B2(new_n387_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n397_), .B2(new_n275_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n392_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n394_), .A2(new_n395_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n393_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT90), .B1(new_n397_), .B2(new_n275_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n385_), .A2(new_n388_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT90), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n310_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n396_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n236_), .A2(new_n275_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n399_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n382_), .B1(new_n401_), .B2(new_n408_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n397_), .A2(KEYINPUT90), .A3(new_n275_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n404_), .B1(new_n403_), .B2(new_n310_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT20), .B(new_n407_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n392_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n413_), .A2(new_n381_), .A3(new_n393_), .A4(new_n400_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n390_), .A2(new_n392_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(new_n412_), .B2(new_n392_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n382_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n414_), .A3(KEYINPUT27), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n338_), .A2(new_n377_), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n361_), .A2(KEYINPUT33), .A3(new_n367_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT94), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n361_), .A2(new_n426_), .A3(KEYINPUT33), .A4(new_n367_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n373_), .B2(new_n366_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n345_), .B(new_n350_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n344_), .A2(new_n346_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n366_), .A3(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n430_), .A2(new_n433_), .A3(new_n414_), .A4(new_n409_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT95), .B1(new_n428_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT33), .B1(new_n361_), .B2(new_n367_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n433_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n415_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT95), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n425_), .A4(new_n427_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n413_), .A2(new_n441_), .A3(new_n393_), .A4(new_n400_), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT96), .Z(new_n443_));
  NAND3_X1  g242(.A1(new_n419_), .A2(KEYINPUT32), .A3(new_n381_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n376_), .A3(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n435_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n332_), .A2(new_n333_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n264_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n423_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G29gat), .B(G36gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G43gat), .B(G50gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G15gat), .B(G22gat), .Z(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT73), .B(G1gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G8gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n459_), .B2(KEYINPUT14), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G1gat), .B(G8gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n454_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n456_), .B1(new_n464_), .B2(new_n455_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT78), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n465_), .A2(new_n468_), .B1(new_n466_), .B2(new_n464_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G169gat), .B(G197gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n469_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G85gat), .B(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT9), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT9), .ZN(new_n479_));
  INV_X1    g278(.A(G92gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n363_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT65), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT6), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT10), .B(G99gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n303_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n478_), .A2(KEYINPUT65), .A3(new_n481_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n486_), .A3(new_n488_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n477_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  OR3_X1    g292(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT7), .ZN(new_n495_));
  OR4_X1    g294(.A1(KEYINPUT66), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n486_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n492_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n493_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n490_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G57gat), .B(G64gat), .Z(new_n501_));
  INV_X1    g300(.A(KEYINPUT11), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n505_));
  XOR2_X1   g304(.A(G71gat), .B(G78gat), .Z(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT68), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n508_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n490_), .B(new_n512_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT64), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n514_), .B(new_n516_), .C1(new_n511_), .C2(new_n510_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  OR2_X1    g317(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n500_), .A2(new_n509_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n518_), .B(new_n520_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G120gat), .B(G148gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G204gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT5), .B(G176gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT13), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n530_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n538_), .A3(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n451_), .A2(new_n476_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n500_), .A2(new_n455_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n454_), .B1(new_n545_), .B2(KEYINPUT72), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT72), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n500_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n550_), .B2(new_n454_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G232gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT34), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(KEYINPUT35), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(KEYINPUT35), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n553_), .A2(KEYINPUT35), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n551_), .B2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n555_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n551_), .A2(new_n562_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n560_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT36), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n566_), .A2(new_n554_), .B1(new_n567_), .B2(new_n558_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT37), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT77), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n509_), .B(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(new_n462_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n462_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT76), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT75), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G183gat), .B(G211gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n572_), .B(new_n462_), .Z(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(KEYINPUT17), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n576_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n582_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n573_), .A2(new_n574_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n591_), .A2(new_n575_), .A3(new_n585_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n570_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n584_), .A2(new_n576_), .A3(new_n586_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n575_), .B1(new_n591_), .B2(new_n585_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(KEYINPUT77), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n558_), .A2(new_n567_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n555_), .B2(new_n563_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n559_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n566_), .A2(new_n600_), .A3(new_n554_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT37), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n569_), .A2(new_n597_), .A3(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n544_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n458_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n376_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT99), .B1(new_n564_), .B2(new_n568_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n599_), .A2(new_n610_), .A3(new_n601_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR4_X1   g412(.A1(new_n451_), .A2(new_n476_), .A3(new_n543_), .A4(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n587_), .A2(new_n592_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n377_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(new_n422_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(new_n615_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n614_), .A2(KEYINPUT100), .A3(new_n615_), .A4(new_n620_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(G8gat), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n623_), .A2(new_n627_), .A3(G8gat), .A4(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(G8gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n605_), .A2(new_n630_), .A3(new_n620_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(KEYINPUT40), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n616_), .B2(new_n449_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n605_), .A2(new_n637_), .A3(new_n449_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n616_), .B2(new_n448_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n605_), .A2(new_n642_), .A3(new_n448_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1327gat));
  NOR2_X1   g445(.A1(new_n612_), .A2(new_n597_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n544_), .A2(new_n647_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n648_), .A2(G29gat), .A3(new_n377_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n597_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n650_), .A2(new_n541_), .A3(new_n475_), .A4(new_n542_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT101), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n446_), .A2(new_n450_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n423_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n569_), .A2(new_n603_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n451_), .A2(KEYINPUT43), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n652_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT44), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(new_n653_), .A3(new_n657_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT43), .B1(new_n451_), .B2(new_n659_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n652_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n376_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(G29gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(G29gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n649_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT103), .B(new_n649_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1328gat));
  NAND3_X1  g475(.A1(new_n663_), .A2(new_n620_), .A3(new_n667_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n648_), .ZN(new_n679_));
  INV_X1    g478(.A(G36gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n620_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n683_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n686_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT46), .B1(new_n686_), .B2(KEYINPUT105), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n648_), .B2(new_n264_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n663_), .A2(G43gat), .A3(new_n449_), .A4(new_n667_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n697_), .B(new_n691_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1330gat));
  NAND3_X1  g500(.A1(new_n663_), .A2(new_n448_), .A3(new_n667_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n663_), .A2(KEYINPUT108), .A3(new_n448_), .A4(new_n667_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(G50gat), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT109), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(G50gat), .A4(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n648_), .A2(G50gat), .A3(new_n447_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1331gat));
  NOR3_X1   g511(.A1(new_n451_), .A2(new_n475_), .A3(new_n650_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n543_), .A3(new_n612_), .ZN(new_n714_));
  INV_X1    g513(.A(G57gat), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n377_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n656_), .A2(KEYINPUT110), .A3(new_n476_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n451_), .B2(new_n475_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n543_), .A3(new_n604_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(new_n377_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n716_), .B1(new_n722_), .B2(new_n715_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n714_), .B2(new_n422_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n422_), .A2(G64gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n721_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n714_), .B2(new_n264_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n449_), .A2(new_n253_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n721_), .B2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n714_), .B2(new_n447_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n448_), .A2(new_n312_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n721_), .B2(new_n734_), .ZN(G1335gat));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n720_), .A2(new_n736_), .A3(new_n543_), .A4(new_n647_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n717_), .A2(new_n719_), .A3(new_n543_), .A4(new_n647_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT111), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n376_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n543_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n475_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n666_), .A2(new_n650_), .A3(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n376_), .A2(G85gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT112), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n741_), .B1(new_n745_), .B2(new_n747_), .ZN(G1336gat));
  NOR3_X1   g547(.A1(new_n744_), .A2(new_n480_), .A3(new_n422_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n740_), .A2(new_n620_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n480_), .ZN(G1337gat));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n449_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n752_), .A2(G99gat), .B1(KEYINPUT114), .B2(KEYINPUT51), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n740_), .A2(new_n487_), .A3(new_n449_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(KEYINPUT113), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n755_), .B(new_n758_), .ZN(G1338gat));
  OAI21_X1  g558(.A(G106gat), .B1(new_n744_), .B2(new_n447_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT52), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(G106gat), .C1(new_n744_), .C2(new_n447_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n447_), .A2(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT115), .B1(new_n740_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  INV_X1    g566(.A(new_n765_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n767_), .B(new_n768_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n764_), .B(new_n772_), .C1(new_n766_), .C2(new_n769_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1339gat));
  OAI21_X1  g573(.A(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n516_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n524_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n524_), .A2(new_n779_), .A3(new_n777_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n524_), .B2(new_n777_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n529_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  INV_X1    g583(.A(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n524_), .A2(new_n779_), .A3(new_n777_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n784_), .B(new_n528_), .C1(new_n787_), .C2(new_n778_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n464_), .A2(new_n467_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n790_));
  MUX2_X1   g589(.A(new_n790_), .B(new_n469_), .S(new_n472_), .Z(new_n791_));
  NAND4_X1  g590(.A1(new_n783_), .A2(new_n530_), .A3(new_n788_), .A4(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n793_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n657_), .A3(new_n795_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n783_), .A2(new_n475_), .A3(new_n788_), .A4(new_n530_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n791_), .A2(new_n536_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n612_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n796_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n615_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  INV_X1    g606(.A(new_n539_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n604_), .A2(new_n807_), .A3(new_n476_), .A4(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n569_), .A2(new_n597_), .A3(new_n476_), .A4(new_n603_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT54), .B1(new_n810_), .B2(new_n539_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n620_), .A2(new_n377_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n337_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT59), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  OAI21_X1  g619(.A(G113gat), .B1(new_n476_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT117), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n612_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n612_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n597_), .B1(new_n827_), .B2(new_n796_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n817_), .C1(new_n828_), .C2(new_n812_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n819_), .A2(new_n821_), .A3(new_n823_), .A4(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n822_), .B1(new_n818_), .B2(new_n476_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT118), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1340gat));
  AND2_X1   g635(.A1(new_n819_), .A2(new_n829_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n543_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  INV_X1    g638(.A(new_n818_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n841_));
  AOI21_X1  g640(.A(G120gat), .B1(new_n543_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT119), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n841_), .B2(G120gat), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n840_), .B(new_n843_), .C1(new_n842_), .C2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n846_), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n840_), .B2(new_n597_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n615_), .A2(G127gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n837_), .B2(new_n849_), .ZN(G1342gat));
  AOI21_X1  g649(.A(G134gat), .B1(new_n840_), .B2(new_n613_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n657_), .A2(G134gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n837_), .B2(new_n852_), .ZN(G1343gat));
  AOI21_X1  g652(.A(new_n812_), .B1(new_n805_), .B2(new_n804_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n854_), .A2(new_n334_), .A3(new_n816_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n475_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n543_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT120), .B(G148gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1345gat));
  NAND2_X1  g659(.A1(new_n855_), .A2(new_n597_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT61), .B(G155gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n855_), .B2(new_n613_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n865_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n659_), .A2(new_n288_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n855_), .B2(new_n868_), .ZN(G1347gat));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n422_), .A2(new_n376_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n264_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n828_), .B2(new_n812_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n448_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n476_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(new_n877_), .B2(new_n203_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n386_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT62), .B(G169gat), .C1(new_n876_), .C2(new_n476_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(G1348gat));
  NAND2_X1  g680(.A1(new_n875_), .A2(new_n543_), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n854_), .A2(new_n220_), .A3(new_n742_), .A4(new_n448_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n882_), .A2(new_n213_), .B1(new_n873_), .B2(new_n883_), .ZN(G1349gat));
  NOR3_X1   g683(.A1(new_n876_), .A2(new_n805_), .A3(new_n229_), .ZN(new_n885_));
  INV_X1    g684(.A(G183gat), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n814_), .A2(new_n447_), .A3(new_n597_), .A4(new_n873_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1350gat));
  NAND3_X1  g687(.A1(new_n875_), .A2(new_n230_), .A3(new_n613_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G190gat), .B1(new_n876_), .B2(new_n659_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1351gat));
  INV_X1    g690(.A(new_n334_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n615_), .B1(new_n827_), .B2(new_n796_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n892_), .B(new_n871_), .C1(new_n893_), .C2(new_n812_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT122), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n334_), .B1(new_n806_), .B2(new_n813_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n871_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n476_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT124), .B1(new_n899_), .B2(G197gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n897_), .B1(new_n896_), .B2(new_n871_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n854_), .A2(KEYINPUT122), .A3(new_n334_), .A4(new_n872_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n475_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  INV_X1    g703(.A(G197gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(G197gat), .B(new_n475_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT123), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n899_), .A2(new_n909_), .A3(G197gat), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n900_), .A2(new_n906_), .B1(new_n908_), .B2(new_n910_), .ZN(G1352gat));
  AOI21_X1  g710(.A(new_n742_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n269_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT125), .B(G204gat), .Z(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n912_), .B2(new_n915_), .ZN(G1353gat));
  AOI21_X1  g715(.A(new_n805_), .B1(new_n895_), .B2(new_n898_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n917_), .B2(new_n918_), .ZN(G1354gat));
  NAND2_X1  g720(.A1(new_n895_), .A2(new_n898_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G218gat), .B1(new_n922_), .B2(new_n613_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n657_), .A2(G218gat), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT126), .Z(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n922_), .B2(new_n925_), .ZN(G1355gat));
endmodule


