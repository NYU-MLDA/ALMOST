//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT10), .B(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n211_), .B2(new_n206_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G85gat), .A3(G92gat), .ZN(new_n214_));
  XOR2_X1   g013(.A(G85gat), .B(G92gat), .Z(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n212_), .B(new_n214_), .C1(new_n213_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NOR3_X1   g017(.A1(KEYINPUT64), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n209_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n207_), .A2(KEYINPUT65), .A3(new_n208_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n218_), .B1(new_n224_), .B2(new_n215_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n209_), .ZN(new_n226_));
  AOI211_X1 g025(.A(KEYINPUT8), .B(new_n216_), .C1(new_n220_), .C2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n217_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n231_));
  XOR2_X1   g030(.A(G71gat), .B(G78gat), .Z(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n231_), .A2(new_n232_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n228_), .A2(new_n236_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n217_), .B(new_n235_), .C1(new_n225_), .C2(new_n227_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT12), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n228_), .A2(new_n240_), .A3(new_n236_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n203_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n237_), .A2(new_n244_), .A3(new_n238_), .ZN(new_n245_));
  OR3_X1    g044(.A1(new_n228_), .A2(new_n244_), .A3(new_n236_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n203_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G120gat), .B(G148gat), .ZN(new_n249_));
  INV_X1    g048(.A(G204gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT5), .B(G176gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n248_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT67), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n254_), .B2(KEYINPUT67), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(KEYINPUT67), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT68), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n259_), .B1(new_n263_), .B2(new_n256_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n202_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n260_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(KEYINPUT13), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT69), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT69), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT26), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT26), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G190gat), .ZN(new_n276_));
  AND2_X1   g075(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n274_), .B(new_n276_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n279_), .A2(new_n282_), .A3(new_n287_), .A4(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT87), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n289_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n297_), .A2(KEYINPUT87), .A3(new_n279_), .A4(new_n287_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n250_), .A2(G197gat), .ZN(new_n300_));
  INV_X1    g099(.A(G197gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G204gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(G211gat), .A2(G218gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G211gat), .A2(G218gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT21), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT85), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n307_), .B1(new_n301_), .B2(G204gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n303_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT21), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n300_), .A2(new_n302_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n302_), .A2(KEYINPUT85), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n312_), .A2(new_n310_), .A3(new_n313_), .A4(KEYINPUT21), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n316_), .A2(KEYINPUT88), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT88), .B1(new_n316_), .B2(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n284_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n295_), .A2(new_n321_), .A3(new_n296_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n322_), .A2(new_n286_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n299_), .A2(new_n315_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT19), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n322_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(G176gat), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G169gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n295_), .A2(new_n321_), .A3(KEYINPUT80), .A4(new_n296_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n273_), .B2(KEYINPUT26), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n275_), .A2(KEYINPUT78), .A3(G190gat), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n336_), .A2(new_n274_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n287_), .A3(new_n297_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n309_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(KEYINPUT89), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT89), .B1(new_n342_), .B2(new_n343_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n325_), .B(new_n329_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n347_), .B(new_n348_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n315_), .B1(new_n299_), .B2(new_n324_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n342_), .B2(new_n343_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n327_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n346_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n355_), .B1(new_n346_), .B2(new_n358_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT27), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n356_), .A2(new_n357_), .A3(new_n327_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n282_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n320_), .A2(new_n323_), .B1(new_n364_), .B2(new_n279_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n328_), .B1(new_n365_), .B2(new_n315_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n327_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n355_), .A2(KEYINPUT91), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n352_), .A2(new_n370_), .A3(new_n354_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n362_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n346_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n327_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n342_), .A2(new_n343_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT89), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n376_), .B1(new_n381_), .B2(new_n366_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT92), .B(new_n372_), .C1(new_n382_), .C2(new_n363_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n374_), .A2(new_n375_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n361_), .B1(new_n384_), .B2(KEYINPUT27), .ZN(new_n385_));
  INV_X1    g184(.A(G141gat), .ZN(new_n386_));
  INV_X1    g185(.A(G148gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G155gat), .ZN(new_n391_));
  INV_X1    g190(.A(G162gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(KEYINPUT83), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(G155gat), .B2(G162gat), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n390_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n393_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT2), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n389_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n403_), .A2(new_n405_), .A3(new_n406_), .A4(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n401_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n401_), .A2(KEYINPUT84), .A3(new_n408_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n400_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT28), .B(G22gat), .ZN(new_n416_));
  INV_X1    g215(.A(G50gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n415_), .B(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G78gat), .B(G106gat), .Z(new_n420_));
  OAI21_X1  g219(.A(new_n343_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n396_), .A2(new_n399_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n390_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n401_), .A2(KEYINPUT84), .A3(new_n408_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT84), .B1(new_n401_), .B2(new_n408_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n315_), .B1(new_n430_), .B2(KEYINPUT29), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n422_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n420_), .B1(new_n424_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n419_), .B1(new_n433_), .B2(KEYINPUT86), .ZN(new_n434_));
  INV_X1    g233(.A(new_n420_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n431_), .A2(new_n422_), .ZN(new_n436_));
  AOI211_X1 g235(.A(new_n423_), .B(new_n315_), .C1(new_n430_), .C2(KEYINPUT29), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n424_), .A2(new_n432_), .A3(new_n420_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n434_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT86), .A4(new_n419_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n342_), .B(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G15gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT81), .B(KEYINPUT30), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n445_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G71gat), .B(G99gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G43gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G127gat), .B(G134gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G120gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n452_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n450_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G29gat), .ZN(new_n459_));
  INV_X1    g258(.A(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT0), .B(G57gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n455_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n430_), .A2(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n455_), .B(new_n427_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(KEYINPUT4), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n430_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n464_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n472_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n478_), .A2(new_n463_), .A3(new_n475_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n458_), .A2(new_n480_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n385_), .A2(new_n443_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n367_), .A2(new_n327_), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n356_), .A2(new_n357_), .A3(new_n327_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n373_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n359_), .B1(new_n486_), .B2(KEYINPUT92), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n483_), .B1(new_n487_), .B2(new_n374_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n480_), .B(new_n443_), .C1(new_n488_), .C2(new_n361_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n463_), .B1(new_n478_), .B2(new_n475_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n359_), .A2(new_n360_), .ZN(new_n493_));
  OAI211_X1 g292(.A(KEYINPUT33), .B(new_n463_), .C1(new_n478_), .C2(new_n475_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n466_), .A2(new_n473_), .A3(new_n467_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n464_), .B(new_n495_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .A4(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n346_), .A2(new_n358_), .A3(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT32), .B(new_n355_), .C1(new_n382_), .C2(new_n363_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n499_), .B(new_n500_), .C1(new_n477_), .C2(new_n479_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n441_), .A2(new_n442_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n489_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n458_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n482_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n228_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n228_), .A2(new_n519_), .B1(new_n511_), .B2(new_n510_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n513_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n520_), .A3(new_n513_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G190gat), .B(G218gat), .Z(new_n525_));
  XOR2_X1   g324(.A(G134gat), .B(G162gat), .Z(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  NAND4_X1  g326(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .A4(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(KEYINPUT36), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT70), .ZN(new_n530_));
  INV_X1    g329(.A(new_n524_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(new_n521_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n522_), .A2(new_n524_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT71), .B1(new_n535_), .B2(new_n530_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT37), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT72), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n538_), .A3(new_n530_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(KEYINPUT72), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .A4(new_n528_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n235_), .B(new_n545_), .Z(new_n546_));
  XOR2_X1   g345(.A(G15gat), .B(G22gat), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT73), .B(G8gat), .Z(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(G1gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT73), .B(G8gat), .ZN(new_n554_));
  INV_X1    g353(.A(G1gat), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n556_), .A2(KEYINPUT74), .A3(new_n549_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n548_), .B1(new_n553_), .B2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G1gat), .B(G8gat), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n551_), .A2(new_n552_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT74), .B1(new_n556_), .B2(new_n549_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n559_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n548_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n546_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G211gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT16), .B(G183gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n568_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n568_), .A2(new_n573_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n507_), .A2(new_n544_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n566_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n517_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT75), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n566_), .B2(new_n516_), .ZN(new_n587_));
  AOI211_X1 g386(.A(KEYINPUT75), .B(new_n517_), .C1(new_n560_), .C2(new_n565_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n585_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT76), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n564_), .B1(new_n563_), .B2(new_n548_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n547_), .B(new_n559_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n516_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n566_), .A2(new_n586_), .A3(new_n516_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT76), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n585_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n583_), .B1(new_n590_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n584_), .A2(new_n519_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n583_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n582_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n596_), .A2(new_n597_), .A3(new_n585_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n597_), .B1(new_n596_), .B2(new_n585_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n603_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n582_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n604_), .A2(new_n610_), .A3(KEYINPUT77), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT77), .B1(new_n604_), .B2(new_n610_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n579_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n272_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT93), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n480_), .B(KEYINPUT94), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n555_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n620_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n265_), .A2(new_n613_), .A3(new_n268_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT95), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n265_), .A2(new_n613_), .A3(new_n625_), .A4(new_n268_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n539_), .A2(new_n540_), .A3(new_n528_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT96), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n629_), .A2(new_n507_), .A3(new_n578_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n624_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n480_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n555_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT97), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n621_), .A2(new_n622_), .A3(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n617_), .A2(new_n554_), .A3(new_n385_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n385_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(G8gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(KEYINPUT98), .B(KEYINPUT39), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n638_), .A2(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n636_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n642_), .B(new_n643_), .Z(G1325gat));
  NAND2_X1  g443(.A1(new_n631_), .A2(new_n458_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G15gat), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT41), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT41), .ZN(new_n648_));
  INV_X1    g447(.A(G15gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n615_), .A2(new_n649_), .A3(new_n458_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n631_), .B2(new_n443_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n615_), .A2(new_n652_), .A3(new_n443_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(G1327gat));
  AND3_X1   g457(.A1(new_n624_), .A2(new_n578_), .A3(new_n626_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n458_), .B1(new_n489_), .B2(new_n504_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(new_n482_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n383_), .A2(new_n375_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n484_), .A2(new_n485_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT92), .B1(new_n664_), .B2(new_n372_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT27), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n361_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n668_), .A2(new_n480_), .A3(new_n503_), .A4(new_n458_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n480_), .A2(new_n442_), .A3(new_n441_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n668_), .A2(new_n670_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT101), .B(new_n669_), .C1(new_n671_), .C2(new_n458_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n662_), .A2(new_n544_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n537_), .A2(new_n676_), .A3(new_n542_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n507_), .A2(KEYINPUT103), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n669_), .B1(new_n671_), .B2(new_n458_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n677_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n678_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n675_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n674_), .B1(new_n673_), .B2(KEYINPUT43), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n659_), .B(KEYINPUT44), .C1(new_n684_), .C2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n624_), .A2(new_n578_), .A3(new_n626_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT103), .B1(new_n507_), .B2(new_n677_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n680_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n543_), .B1(new_n680_), .B2(new_n660_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n676_), .B1(new_n691_), .B2(new_n672_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(new_n674_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n685_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n687_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n686_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(G29gat), .A3(new_n618_), .ZN(new_n700_));
  INV_X1    g499(.A(G29gat), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n507_), .A2(new_n627_), .A3(new_n577_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n269_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n613_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n704_), .B2(new_n480_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1328gat));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n385_), .B(new_n686_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT106), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n713_), .A3(G36gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n704_), .A2(G36gat), .A3(new_n668_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n717_));
  XOR2_X1   g516(.A(new_n716_), .B(new_n717_), .Z(new_n718_));
  AOI21_X1  g517(.A(new_n709_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n710_), .A2(new_n713_), .A3(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n713_), .B1(new_n710_), .B2(G36gat), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n718_), .B(new_n709_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n719_), .A2(new_n723_), .ZN(G1329gat));
  NOR3_X1   g523(.A1(new_n704_), .A2(G43gat), .A3(new_n506_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n699_), .A2(new_n458_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G43gat), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1330gat));
  OAI21_X1  g528(.A(G50gat), .B1(new_n698_), .B2(new_n503_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n443_), .A2(new_n417_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n704_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT110), .ZN(G1331gat));
  INV_X1    g532(.A(new_n272_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n613_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n630_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n480_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n703_), .A2(new_n613_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n579_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n618_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT111), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n385_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G64gat), .B1(new_n736_), .B2(new_n668_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT48), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT48), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n750_), .A3(new_n458_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G71gat), .B1(new_n736_), .B2(new_n506_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT49), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT49), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n739_), .A2(new_n756_), .A3(new_n443_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G78gat), .B1(new_n736_), .B2(new_n503_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(KEYINPUT50), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(KEYINPUT50), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1335gat));
  NAND2_X1  g560(.A1(new_n735_), .A2(new_n702_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G85gat), .B1(new_n763_), .B2(new_n618_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n693_), .A2(new_n694_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n578_), .A3(new_n738_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n480_), .A2(new_n460_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  AOI21_X1  g568(.A(G92gat), .B1(new_n763_), .B2(new_n385_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n385_), .A2(G92gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n767_), .B2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n766_), .B2(new_n506_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n458_), .A2(new_n211_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n762_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g575(.A1(new_n503_), .A2(G106gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OR3_X1    g577(.A1(new_n762_), .A2(KEYINPUT112), .A3(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n762_), .B2(new_n778_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G106gat), .B1(new_n766_), .B2(new_n503_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(KEYINPUT52), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT52), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n781_), .B(new_n787_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  NOR3_X1   g588(.A1(new_n613_), .A2(new_n544_), .A3(new_n578_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n703_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n237_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n247_), .B1(new_n794_), .B2(new_n241_), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n795_), .A2(KEYINPUT113), .A3(KEYINPUT55), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT113), .B1(new_n795_), .B2(KEYINPUT55), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n794_), .A2(KEYINPUT114), .A3(new_n241_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n247_), .A3(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .A4(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n253_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n613_), .A2(new_n809_), .A3(new_n254_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n583_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n601_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n596_), .A2(KEYINPUT115), .A3(new_n600_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n602_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n815_), .A3(new_n582_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n610_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT116), .B1(new_n816_), .B2(new_n610_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n819_), .A2(new_n820_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n810_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n822_), .B2(new_n627_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n819_), .A2(new_n820_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n254_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n807_), .A2(KEYINPUT117), .A3(new_n808_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n808_), .A2(KEYINPUT117), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n827_), .A2(KEYINPUT58), .A3(new_n828_), .A4(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n829_), .B(new_n254_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n828_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(new_n544_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  INV_X1    g635(.A(new_n627_), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n836_), .B(new_n837_), .C1(new_n810_), .C2(new_n821_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n824_), .A2(new_n835_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n793_), .B1(new_n840_), .B2(new_n578_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n385_), .A2(new_n443_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n458_), .A3(new_n618_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n613_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n843_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n613_), .A2(G113gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n849_), .B2(new_n850_), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n272_), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G120gat), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(KEYINPUT60), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n703_), .B2(KEYINPUT60), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(KEYINPUT118), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n844_), .B(new_n857_), .C1(KEYINPUT118), .C2(new_n856_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n844_), .B2(new_n577_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n577_), .A2(G127gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n849_), .B2(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n844_), .B2(new_n629_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n544_), .A2(G134gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n849_), .B2(new_n864_), .ZN(G1343gat));
  NAND3_X1  g664(.A1(new_n618_), .A2(new_n443_), .A3(new_n506_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n841_), .A2(new_n385_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n613_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n272_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(G148gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1345gat));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n577_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  AOI21_X1  g674(.A(G162gat), .B1(new_n867_), .B2(new_n629_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n543_), .A2(new_n392_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n867_), .B2(new_n877_), .ZN(G1347gat));
  NOR3_X1   g677(.A1(new_n618_), .A2(new_n668_), .A3(new_n506_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n880_), .A2(KEYINPUT120), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT120), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n503_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n823_), .A2(new_n838_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n577_), .B1(new_n885_), .B2(new_n835_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n613_), .B(new_n884_), .C1(new_n886_), .C2(new_n793_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n283_), .B1(new_n887_), .B2(KEYINPUT121), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n840_), .A2(new_n578_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n793_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(new_n613_), .A4(new_n884_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n888_), .A2(new_n889_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n889_), .B1(new_n888_), .B2(new_n894_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(KEYINPUT122), .A3(new_n884_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n841_), .B2(new_n883_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n613_), .B1(new_n319_), .B2(new_n318_), .ZN(new_n901_));
  OAI22_X1  g700(.A1(new_n895_), .A2(new_n896_), .B1(new_n900_), .B2(new_n901_), .ZN(G1348gat));
  NOR4_X1   g701(.A1(new_n841_), .A2(new_n284_), .A3(new_n734_), .A4(new_n883_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n897_), .A2(new_n269_), .A3(new_n899_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n284_), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n578_), .A2(new_n336_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n897_), .A2(new_n899_), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n577_), .B(new_n884_), .C1(new_n886_), .C2(new_n793_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G183gat), .B1(new_n910_), .B2(KEYINPUT124), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(KEYINPUT124), .B2(new_n910_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n897_), .A2(new_n899_), .A3(KEYINPUT123), .A4(new_n906_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n909_), .A2(new_n912_), .A3(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n900_), .B2(new_n543_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n629_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT125), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n900_), .B2(new_n917_), .ZN(G1351gat));
  AND3_X1   g717(.A1(new_n385_), .A2(new_n670_), .A3(new_n506_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n892_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n613_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  OAI211_X1 g721(.A(new_n920_), .B(new_n272_), .C1(KEYINPUT126), .C2(new_n250_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n920_), .A2(new_n272_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT126), .B(G204gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(G1353gat));
  NAND2_X1  g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n920_), .A2(new_n577_), .A3(new_n927_), .ZN(new_n928_));
  OR2_X1    g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1354gat));
  NAND3_X1  g729(.A1(new_n892_), .A2(new_n629_), .A3(new_n919_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n932_));
  AOI21_X1  g731(.A(G218gat), .B1(new_n931_), .B2(KEYINPUT127), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n544_), .A2(G218gat), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n932_), .A2(new_n933_), .B1(new_n920_), .B2(new_n934_), .ZN(G1355gat));
endmodule


