//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n979_, new_n980_, new_n982_, new_n983_, new_n984_, new_n986_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n992_, new_n994_,
    new_n995_;
  INV_X1    g000(.A(KEYINPUT108), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT23), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n217_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n218_), .C2(new_n219_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n222_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n218_), .A2(new_n219_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n213_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G169gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n212_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT95), .ZN(new_n237_));
  XOR2_X1   g036(.A(G211gat), .B(G218gat), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G204gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(G197gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT90), .B(G204gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n242_), .B2(G197gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT92), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(G197gat), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n241_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n248_), .A2(KEYINPUT92), .A3(new_n244_), .A4(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n239_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G197gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G197gat), .A2(G204gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT21), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n254_), .A2(KEYINPUT91), .A3(KEYINPUT21), .A4(new_n255_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT93), .B1(new_n252_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n248_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT92), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n238_), .B1(new_n264_), .B2(new_n250_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT93), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n259_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n243_), .A2(KEYINPUT94), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n248_), .A2(new_n249_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT94), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n270_), .A2(new_n273_), .A3(KEYINPUT21), .A4(new_n238_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n237_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT95), .B(new_n276_), .C1(new_n261_), .C2(new_n268_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n227_), .B(new_n236_), .C1(new_n275_), .C2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n274_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n218_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT25), .B1(new_n218_), .B2(KEYINPUT80), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n224_), .A2(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n231_), .B(new_n217_), .C1(new_n283_), .C2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT22), .B1(new_n211_), .B2(KEYINPUT82), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT82), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT22), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(G169gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n290_), .A3(new_n212_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n213_), .B1(new_n291_), .B2(KEYINPUT83), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n223_), .A2(new_n232_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n287_), .A2(new_n290_), .A3(new_n294_), .A4(new_n212_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n286_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n279_), .B1(new_n282_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n210_), .B1(new_n278_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n233_), .A2(KEYINPUT98), .A3(new_n235_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT98), .B1(new_n233_), .B2(new_n235_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n227_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n282_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n298_), .A2(new_n299_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n269_), .A2(new_n308_), .A3(new_n274_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT20), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n209_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n207_), .B1(new_n302_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n276_), .B1(new_n261_), .B2(new_n268_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n227_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n305_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n303_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n301_), .A2(new_n210_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n207_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT99), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n310_), .A2(new_n320_), .A3(new_n209_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n310_), .B2(new_n209_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n318_), .B(new_n319_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n312_), .A2(new_n323_), .A3(KEYINPUT27), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT101), .ZN(new_n326_));
  INV_X1    g125(.A(new_n318_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n313_), .B2(new_n316_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n282_), .A2(new_n300_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n209_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT99), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n310_), .A2(new_n320_), .A3(new_n209_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n326_), .B1(new_n333_), .B2(new_n319_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n318_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT101), .A3(new_n207_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n336_), .A3(new_n323_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n325_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G50gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT89), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(KEYINPUT86), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT86), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(G141gat), .A3(G148gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n351_), .B2(new_n346_), .ZN(new_n352_));
  INV_X1    g151(.A(G141gat), .ZN(new_n353_));
  INV_X1    g152(.A(G148gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT87), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT87), .A4(KEYINPUT3), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n352_), .A2(KEYINPUT88), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT88), .B1(new_n352_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n344_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n342_), .A2(KEYINPUT1), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n342_), .A2(KEYINPUT1), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n341_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n353_), .A2(new_n354_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n351_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT28), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n369_));
  INV_X1    g168(.A(G22gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n362_), .A2(new_n371_), .A3(new_n372_), .A4(new_n367_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n370_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n370_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n340_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(G50gat), .A3(new_n374_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT97), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n282_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n282_), .A2(KEYINPUT95), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n269_), .A2(new_n237_), .A3(new_n274_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n368_), .A2(KEYINPUT29), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n384_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n390_), .B2(new_n384_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n386_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n382_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n377_), .A2(new_n379_), .A3(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n383_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n383_), .B2(new_n396_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n202_), .B1(new_n339_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G127gat), .B(G134gat), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n402_), .A2(G113gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(G113gat), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n403_), .A2(G120gat), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(G120gat), .B1(new_n403_), .B2(new_n404_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n343_), .B(KEYINPUT89), .Z(new_n408_));
  AOI21_X1  g207(.A(new_n349_), .B1(G141gat), .B2(G148gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n345_), .A2(KEYINPUT86), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n346_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n347_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n359_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n352_), .A2(KEYINPUT88), .A3(new_n359_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n408_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n367_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n407_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n405_), .A2(new_n406_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n362_), .A2(new_n420_), .A3(new_n367_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(KEYINPUT4), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT102), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n419_), .A2(KEYINPUT4), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT102), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n419_), .A2(new_n421_), .A3(new_n425_), .A4(KEYINPUT4), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n419_), .A2(new_n421_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT103), .B(G85gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT0), .B(G57gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT106), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n432_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n439_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n434_), .A2(new_n441_), .A3(new_n439_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n308_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT30), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(KEYINPUT85), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(KEYINPUT85), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n420_), .B(KEYINPUT31), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n456_), .A2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n339_), .A2(new_n399_), .A3(new_n202_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n401_), .A2(new_n447_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n431_), .B(KEYINPUT104), .Z(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n429_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n443_), .C1(new_n429_), .C2(new_n427_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n334_), .A2(new_n336_), .A3(new_n466_), .A4(new_n323_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n440_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n311_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n301_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n314_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n236_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n470_), .B1(new_n473_), .B2(new_n210_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT105), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT105), .B(new_n476_), .C1(new_n302_), .C2(new_n311_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n333_), .A2(new_n475_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n445_), .A2(new_n446_), .A3(new_n481_), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n467_), .A2(new_n469_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT107), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n399_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n483_), .B2(new_n399_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n397_), .A2(new_n398_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n339_), .A2(new_n447_), .A3(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n485_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n463_), .B1(new_n489_), .B2(new_n461_), .ZN(new_n490_));
  AND2_X1   g289(.A1(G57gat), .A2(G64gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G57gat), .A2(G64gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT11), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT68), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT68), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(KEYINPUT11), .C1(new_n491_), .C2(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n494_), .ZN(new_n499_));
  INV_X1    g298(.A(G71gat), .ZN(new_n500_));
  INV_X1    g299(.A(G78gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n493_), .A2(new_n494_), .B1(G71gat), .B2(G78gat), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(new_n495_), .A3(new_n502_), .A4(new_n497_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT10), .B(G99gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT64), .B(G106gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT66), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT65), .B(G85gat), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G92gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G92gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G85gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G92gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n515_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT9), .ZN(new_n527_));
  OR2_X1    g326(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n528_), .A2(new_n517_), .A3(G92gat), .A4(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(KEYINPUT66), .A3(new_n530_), .ZN(new_n531_));
  AOI211_X1 g330(.A(new_n511_), .B(new_n514_), .C1(new_n525_), .C2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n533_));
  NOR2_X1   g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n526_), .B(new_n533_), .C1(new_n511_), .C2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n509_), .B(KEYINPUT6), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(new_n537_), .A3(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n540_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n526_), .A3(new_n533_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n508_), .B1(new_n532_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n514_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n531_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT66), .B1(new_n527_), .B2(new_n530_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n542_), .B(new_n548_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n505_), .A2(new_n507_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n541_), .A4(new_n545_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n553_), .A3(KEYINPUT12), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n551_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n508_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G230gat), .A2(G233gat), .ZN(new_n560_));
  MUX2_X1   g359(.A(new_n554_), .B(new_n559_), .S(new_n560_), .Z(new_n561_));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G176gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n240_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n565_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(KEYINPUT69), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT69), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n561_), .A2(new_n569_), .A3(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(KEYINPUT13), .A3(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G29gat), .B(G36gat), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G43gat), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n580_), .B(KEYINPUT71), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(G43gat), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n340_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(G43gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(new_n583_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(G50gat), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592_));
  INV_X1    g391(.A(G1gat), .ZN(new_n593_));
  INV_X1    g392(.A(G8gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT14), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G1gat), .B(G8gat), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n596_), .B(new_n597_), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n587_), .A2(new_n590_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(KEYINPUT78), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT78), .B1(new_n599_), .B2(new_n602_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n579_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n600_), .A2(new_n601_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT15), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n587_), .A2(KEYINPUT15), .A3(new_n590_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n607_), .B1(new_n611_), .B2(new_n601_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n578_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n577_), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n577_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n211_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n253_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n614_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n612_), .A2(new_n578_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT78), .ZN(new_n623_));
  INV_X1    g422(.A(new_n602_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(new_n607_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n578_), .B1(new_n625_), .B2(new_n603_), .ZN(new_n626_));
  OAI21_X1  g425(.A(KEYINPUT79), .B1(new_n622_), .B2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n621_), .B1(new_n627_), .B2(new_n615_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n620_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n576_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G190gat), .B(G218gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT70), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT34), .ZN(new_n636_));
  INV_X1    g435(.A(new_n556_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n600_), .A2(new_n556_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT35), .B(new_n636_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n610_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT15), .B1(new_n587_), .B2(new_n590_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n556_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n636_), .A2(KEYINPUT35), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n636_), .A2(KEYINPUT35), .ZN(new_n645_));
  INV_X1    g444(.A(new_n639_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .A4(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT36), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n633_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n649_), .A3(new_n633_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n652_), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT36), .B(new_n632_), .C1(new_n640_), .C2(new_n647_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n650_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n640_), .A2(new_n647_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(KEYINPUT37), .A3(new_n660_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n598_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(new_n552_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT75), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT17), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(G183gat), .B(G211gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(G127gat), .B(G155gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n674_), .B(new_n675_), .Z(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT74), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n668_), .A2(new_n679_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n680_), .A2(new_n670_), .A3(KEYINPUT17), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n669_), .A2(new_n670_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n680_), .A2(KEYINPUT17), .A3(new_n676_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n678_), .A2(new_n681_), .A3(new_n682_), .A4(new_n683_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n684_), .A2(KEYINPUT76), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(KEYINPUT76), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(KEYINPUT77), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT77), .B1(new_n685_), .B2(new_n686_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n665_), .A2(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n490_), .A2(new_n631_), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n447_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n593_), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT38), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n483_), .A2(new_n399_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT107), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n339_), .A2(new_n447_), .A3(new_n487_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n483_), .A2(new_n484_), .A3(new_n399_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n339_), .A2(new_n399_), .A3(new_n202_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(new_n400_), .A3(new_n460_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n460_), .A2(new_n701_), .B1(new_n703_), .B2(new_n447_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n696_), .B1(new_n704_), .B2(new_n661_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n661_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n490_), .A2(KEYINPUT109), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n685_), .A2(new_n686_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n631_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G1gat), .B1(new_n710_), .B2(new_n447_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n695_), .A2(new_n711_), .ZN(G1324gat));
  INV_X1    g511(.A(new_n339_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n692_), .A2(new_n594_), .A3(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n708_), .A2(new_n709_), .A3(new_n713_), .A4(new_n631_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT39), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(G8gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G8gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT40), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT40), .B(new_n714_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1325gat));
  INV_X1    g522(.A(G15gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n692_), .A2(new_n724_), .A3(new_n461_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n710_), .A2(new_n460_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT41), .B1(new_n726_), .B2(G15gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1326gat));
  NAND2_X1  g528(.A1(new_n487_), .A2(new_n370_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT110), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n692_), .A2(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n710_), .A2(new_n399_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(G22gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n733_), .B2(G22gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1327gat));
  INV_X1    g536(.A(G29gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n663_), .A2(new_n664_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n704_), .B2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n490_), .A2(KEYINPUT43), .A3(new_n665_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(new_n631_), .A3(new_n742_), .A4(new_n690_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT44), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n738_), .B1(new_n744_), .B2(new_n693_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n689_), .A2(new_n706_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n490_), .A2(new_n631_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n490_), .A2(KEYINPUT111), .A3(new_n631_), .A4(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n751_), .A2(G29gat), .A3(new_n447_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n745_), .A2(new_n752_), .ZN(G1328gat));
  NAND2_X1  g552(.A1(new_n701_), .A2(new_n460_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n739_), .B(new_n740_), .C1(new_n754_), .C2(new_n463_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT43), .B1(new_n490_), .B2(new_n665_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n757_), .A2(KEYINPUT44), .A3(new_n631_), .A4(new_n690_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n743_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n758_), .A2(new_n713_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G36gat), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n339_), .A2(G36gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n749_), .A2(new_n750_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT112), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n749_), .A2(new_n766_), .A3(new_n750_), .A4(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(KEYINPUT45), .A3(new_n767_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n762_), .A2(new_n770_), .A3(KEYINPUT46), .A4(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1329gat));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n758_), .A2(new_n461_), .A3(new_n760_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G43gat), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n461_), .A2(new_n583_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n751_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n779_), .B(KEYINPUT47), .C1(new_n751_), .C2(new_n781_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1330gat));
  NAND2_X1  g584(.A1(new_n744_), .A2(new_n487_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n744_), .A2(new_n788_), .A3(new_n487_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(G50gat), .A3(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n749_), .A2(new_n340_), .A3(new_n487_), .A4(new_n750_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1331gat));
  NOR2_X1   g591(.A1(new_n575_), .A2(new_n629_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n704_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n691_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G57gat), .B1(new_n797_), .B2(new_n693_), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n690_), .B(new_n794_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n693_), .A2(G57gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(G1332gat));
  INV_X1    g600(.A(G64gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n802_), .A3(new_n713_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT48), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(new_n713_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G64gat), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT48), .B(new_n802_), .C1(new_n799_), .C2(new_n713_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(G1333gat));
  NAND3_X1  g607(.A1(new_n797_), .A2(new_n500_), .A3(new_n461_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n799_), .A2(new_n461_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(G71gat), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT49), .B(new_n500_), .C1(new_n799_), .C2(new_n461_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(G1334gat));
  NAND3_X1  g613(.A1(new_n797_), .A2(new_n501_), .A3(new_n487_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n799_), .A2(new_n487_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G78gat), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(KEYINPUT50), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(KEYINPUT50), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n815_), .B1(new_n818_), .B2(new_n819_), .ZN(G1335gat));
  NAND4_X1  g619(.A1(new_n741_), .A2(new_n690_), .A3(new_n742_), .A4(new_n793_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n821_), .A2(new_n447_), .A3(new_n516_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT114), .B1(new_n795_), .B2(new_n746_), .ZN(new_n823_));
  AND4_X1   g622(.A1(KEYINPUT114), .A2(new_n490_), .A3(new_n746_), .A4(new_n793_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n693_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n826_), .B2(new_n522_), .ZN(G1336gat));
  NOR3_X1   g626(.A1(new_n821_), .A2(new_n520_), .A3(new_n339_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n713_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n520_), .ZN(G1337gat));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n461_), .A3(new_n512_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G99gat), .B1(new_n821_), .B2(new_n460_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g633(.A(G106gat), .B1(new_n821_), .B2(new_n399_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n836_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n487_), .B(new_n513_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT115), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n840_), .B(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n837_), .A4(new_n838_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1339gat));
  INV_X1    g646(.A(new_n560_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n555_), .A2(new_n848_), .A3(new_n558_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n555_), .A2(KEYINPUT116), .A3(new_n558_), .A4(new_n848_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT55), .B(new_n848_), .C1(new_n555_), .C2(new_n558_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n851_), .A2(new_n853_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n849_), .A2(new_n850_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n852_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n861_), .B(KEYINPUT117), .C1(new_n855_), .C2(new_n856_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n565_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n863_), .A2(new_n866_), .A3(new_n864_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n865_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n620_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n578_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n612_), .A2(new_n579_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n619_), .A3(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n566_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n869_), .A2(KEYINPUT58), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n863_), .A2(new_n864_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n868_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n863_), .A2(new_n866_), .A3(new_n864_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n879_), .B1(new_n883_), .B2(new_n874_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n869_), .A2(KEYINPUT120), .A3(new_n875_), .A4(KEYINPUT58), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n878_), .A2(new_n665_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT121), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n740_), .B1(new_n877_), .B2(new_n876_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n566_), .B1(new_n620_), .B2(new_n628_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n863_), .A2(new_n864_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n865_), .ZN(new_n893_));
  AND4_X1   g692(.A1(new_n870_), .A2(new_n570_), .A3(new_n568_), .A4(new_n873_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n706_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  OR2_X1    g694(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n887_), .A2(new_n890_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n709_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n740_), .A2(new_n630_), .A3(new_n689_), .A4(new_n575_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n904_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n703_), .A2(new_n693_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G113gat), .B1(new_n908_), .B2(new_n629_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(KEYINPUT59), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n897_), .A2(new_n886_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n690_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT122), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n914_), .A3(new_n690_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n904_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(new_n917_), .A3(new_n906_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n910_), .A2(new_n918_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n629_), .A2(G113gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n909_), .B1(new_n919_), .B2(new_n920_), .ZN(G1340gat));
  NAND3_X1  g720(.A1(new_n910_), .A2(new_n918_), .A3(new_n576_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT123), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n910_), .A2(new_n918_), .A3(new_n924_), .A4(new_n576_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(G120gat), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(G120gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n908_), .B(new_n928_), .C1(KEYINPUT60), .C2(new_n927_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n929_), .ZN(G1341gat));
  AOI21_X1  g729(.A(G127gat), .B1(new_n908_), .B2(new_n689_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n709_), .A2(G127gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n919_), .B2(new_n932_), .ZN(G1342gat));
  NAND3_X1  g732(.A1(new_n919_), .A2(G134gat), .A3(new_n665_), .ZN(new_n934_));
  INV_X1    g733(.A(G134gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n907_), .B2(new_n706_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n937_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n934_), .A2(new_n938_), .A3(new_n939_), .ZN(G1343gat));
  AOI21_X1  g739(.A(new_n903_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n461_), .ZN(new_n942_));
  AND4_X1   g741(.A1(new_n693_), .A2(new_n942_), .A3(new_n487_), .A4(new_n339_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n629_), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT125), .B(G141gat), .Z(new_n945_));
  XNOR2_X1  g744(.A(new_n944_), .B(new_n945_), .ZN(G1344gat));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n576_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g747(.A1(new_n943_), .A2(new_n689_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT61), .B(G155gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1346gat));
  AOI21_X1  g750(.A(G162gat), .B1(new_n943_), .B2(new_n661_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n665_), .A2(G162gat), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n943_), .B2(new_n953_), .ZN(G1347gat));
  NOR3_X1   g753(.A1(new_n339_), .A2(new_n693_), .A3(new_n460_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n916_), .A2(new_n399_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n211_), .B1(new_n956_), .B2(new_n629_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n916_), .A2(new_n399_), .A3(new_n955_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n234_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n958_), .A2(new_n959_), .A3(new_n630_), .ZN(new_n960_));
  OAI21_X1  g759(.A(KEYINPUT62), .B1(new_n957_), .B2(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(KEYINPUT62), .B2(new_n957_), .ZN(G1348gat));
  AOI21_X1  g761(.A(G176gat), .B1(new_n956_), .B2(new_n576_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n905_), .A2(new_n964_), .A3(new_n399_), .ZN(new_n965_));
  OAI21_X1  g764(.A(KEYINPUT126), .B1(new_n941_), .B2(new_n487_), .ZN(new_n966_));
  AND3_X1   g765(.A1(new_n965_), .A2(new_n955_), .A3(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n575_), .A2(new_n212_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n963_), .B1(new_n967_), .B2(new_n968_), .ZN(G1349gat));
  NAND4_X1  g768(.A1(new_n965_), .A2(new_n966_), .A3(new_n689_), .A4(new_n955_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n218_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n225_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n956_), .A2(new_n709_), .A3(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n971_), .A2(new_n973_), .A3(new_n976_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n977_), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n956_), .A2(new_n224_), .A3(new_n661_), .ZN(new_n979_));
  OAI21_X1  g778(.A(G190gat), .B1(new_n958_), .B2(new_n740_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1351gat));
  NOR2_X1   g780(.A1(new_n339_), .A2(new_n693_), .ZN(new_n982_));
  AND3_X1   g781(.A1(new_n942_), .A2(new_n487_), .A3(new_n982_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(new_n629_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g784(.A1(new_n983_), .A2(new_n576_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(new_n242_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n987_), .B1(new_n986_), .B2(new_n240_), .ZN(G1353gat));
  NAND2_X1  g787(.A1(new_n983_), .A2(new_n709_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(KEYINPUT63), .B(G211gat), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n989_), .A2(new_n990_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n991_), .B1(new_n989_), .B2(new_n992_), .ZN(G1354gat));
  AOI21_X1  g792(.A(G218gat), .B1(new_n983_), .B2(new_n661_), .ZN(new_n994_));
  AND2_X1   g793(.A1(new_n665_), .A2(G218gat), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n994_), .B1(new_n983_), .B2(new_n995_), .ZN(G1355gat));
endmodule


