// Benchmark "c7552" written by ABC on Wed Jul  6 02:19:16 2022

module c7552 ( 
    G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47,
    G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65,
    G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83,
    G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110,
    G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134,
    G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156,
    G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168,
    G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216,
    G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228,
    G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240,
    G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496,
    G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253,
    G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743,
    G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432,
    G4437, G4526, G4528,
    G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399  );
  input  G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41,
    G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63,
    G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81,
    G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106,
    G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130,
    G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154,
    G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166,
    G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190,
    G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202,
    G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214,
    G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226,
    G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238,
    G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486,
    G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239,
    G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729,
    G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420,
    G4427, G4432, G4437, G4526, G4528;
  output G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490,
    G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550,
    G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524,
    G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284,
    G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270,
    G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249,
    G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336,
    G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359,
    G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399;
  wire new_n362_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1033_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1332_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1357_,
    new_n1359_, new_n1360_, new_n1361_, new_n1363_, new_n1364_, new_n1365_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1389_, new_n1391_, new_n1392_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1424_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_;
  BUF_X1    g0000(.A(G1), .Z(G2));
  BUF_X1    g0001(.A(G1), .Z(G3));
  BUF_X1    g0002(.A(G1459), .Z(G450));
  BUF_X1    g0003(.A(G1469), .Z(G448));
  BUF_X1    g0004(.A(G1480), .Z(G444));
  BUF_X1    g0005(.A(G1486), .Z(G442));
  BUF_X1    g0006(.A(G1492), .Z(G440));
  BUF_X1    g0007(.A(G1496), .Z(G438));
  BUF_X1    g0008(.A(G2208), .Z(G496));
  BUF_X1    g0009(.A(G2218), .Z(G494));
  BUF_X1    g0010(.A(G2224), .Z(G492));
  BUF_X1    g0011(.A(G2230), .Z(G490));
  BUF_X1    g0012(.A(G2236), .Z(G488));
  BUF_X1    g0013(.A(G2239), .Z(G486));
  BUF_X1    g0014(.A(G2247), .Z(G484));
  BUF_X1    g0015(.A(G2253), .Z(G482));
  BUF_X1    g0016(.A(G2256), .Z(G480));
  BUF_X1    g0017(.A(G3698), .Z(G560));
  BUF_X1    g0018(.A(G3701), .Z(G542));
  BUF_X1    g0019(.A(G3705), .Z(G558));
  BUF_X1    g0020(.A(G3711), .Z(G556));
  BUF_X1    g0021(.A(G3717), .Z(G554));
  BUF_X1    g0022(.A(G3723), .Z(G552));
  BUF_X1    g0023(.A(G3729), .Z(G550));
  BUF_X1    g0024(.A(G3737), .Z(G548));
  BUF_X1    g0025(.A(G3743), .Z(G546));
  BUF_X1    g0026(.A(G3749), .Z(G544));
  BUF_X1    g0027(.A(G4393), .Z(G540));
  BUF_X1    g0028(.A(G4400), .Z(G538));
  BUF_X1    g0029(.A(G4405), .Z(G536));
  BUF_X1    g0030(.A(G4410), .Z(G534));
  BUF_X1    g0031(.A(G4415), .Z(G532));
  BUF_X1    g0032(.A(G4420), .Z(G530));
  BUF_X1    g0033(.A(G4427), .Z(G528));
  BUF_X1    g0034(.A(G4432), .Z(G526));
  BUF_X1    g0035(.A(G4437), .Z(G524));
  INV_X1    g0036(.A(G15), .ZN(G279));
  BUF_X1    g0037(.A(G1462), .Z(G436));
  BUF_X1    g0038(.A(G2211), .Z(G478));
  BUF_X1    g0039(.A(G4394), .Z(G522));
  OR2_X1    g0040(.A1(G5), .A2(G57), .ZN(G402));
  NAND4_X1  g0041(.A1(G150), .A2(G184), .A3(G228), .A4(G240), .ZN(G404));
  NAND4_X1  g0042(.A1(G152), .A2(G210), .A3(G218), .A4(G230), .ZN(G406));
  NAND4_X1  g0043(.A1(G182), .A2(G183), .A3(G185), .A4(G186), .ZN(G408));
  NAND4_X1  g0044(.A1(G162), .A2(G172), .A3(G188), .A4(G199), .ZN(G410));
  BUF_X1    g0045(.A(G1), .Z(G432));
  BUF_X1    g0046(.A(G106), .Z(G446));
  INV_X1    g0047(.A(G5), .ZN(new_n362_));
  NAND2_X1  g0048(.A1(new_n362_), .A2(G1197), .ZN(G284));
  INV_X1    g0049(.A(G15), .ZN(G286));
  NAND2_X1  g0050(.A1(new_n362_), .A2(G1197), .ZN(G289));
  NAND3_X1  g0051(.A1(new_n362_), .A2(G133), .A3(G134), .ZN(G292));
  INV_X1    g0052(.A(G15), .ZN(G341));
  NAND3_X1  g0053(.A1(new_n362_), .A2(G133), .A3(G134), .ZN(G281));
  BUF_X1    g0054(.A(G1), .Z(G453));
  AND2_X1   g0055(.A1(G1), .A2(G163), .ZN(G278));
  INV_X1    g0056(.A(G18), .ZN(new_n371_));
  NAND2_X1  g0057(.A1(new_n371_), .A2(G41), .ZN(new_n372_));
  NAND2_X1  g0058(.A1(new_n371_), .A2(G3701), .ZN(new_n373_));
  XNOR2_X1  g0059(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g0060(.A(G4526), .ZN(new_n375_));
  XNOR2_X1  g0061(.A(new_n374_), .B(new_n375_), .ZN(G373));
  AND2_X1   g0062(.A1(G9), .A2(G12), .ZN(new_n377_));
  INV_X1    g0063(.A(G213), .ZN(new_n378_));
  AOI21_X1  g0064(.A(new_n377_), .B1(G18), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g0065(.A(G1486), .ZN(new_n380_));
  XNOR2_X1  g0066(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g0067(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g0068(.A1(G9), .A2(G12), .ZN(new_n383_));
  OAI21_X1  g0069(.A(new_n383_), .B1(new_n371_), .B2(G215), .ZN(new_n384_));
  INV_X1    g0070(.A(G106), .ZN(new_n385_));
  NAND2_X1  g0071(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g0072(.A(new_n383_), .B(G106), .C1(new_n371_), .C2(G215), .ZN(new_n387_));
  NAND2_X1  g0073(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g0074(.A(new_n383_), .B1(new_n371_), .B2(G216), .ZN(new_n389_));
  INV_X1    g0075(.A(G1469), .ZN(new_n390_));
  NAND2_X1  g0076(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g0077(.A(new_n383_), .B(G1469), .C1(new_n371_), .C2(G216), .ZN(new_n392_));
  NAND2_X1  g0078(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g0079(.A1(new_n382_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g0080(.A(new_n383_), .B1(new_n371_), .B2(G209), .ZN(new_n395_));
  INV_X1    g0081(.A(G1462), .ZN(new_n396_));
  XNOR2_X1  g0082(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g0083(.A(new_n397_), .ZN(new_n398_));
  OAI21_X1  g0084(.A(new_n383_), .B1(new_n371_), .B2(G214), .ZN(new_n399_));
  INV_X1    g0085(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g0086(.A1(new_n400_), .A2(G1480), .ZN(new_n401_));
  INV_X1    g0087(.A(G1480), .ZN(new_n402_));
  NAND2_X1  g0088(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g0089(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g0090(.A(new_n404_), .ZN(new_n405_));
  NOR3_X1   g0091(.A1(new_n394_), .A2(new_n398_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g0092(.A1(G1492), .A2(G4528), .ZN(new_n407_));
  XNOR2_X1  g0093(.A(new_n407_), .B(G38), .ZN(new_n408_));
  NAND2_X1  g0094(.A1(G1496), .A2(G4528), .ZN(new_n409_));
  XNOR2_X1  g0095(.A(new_n409_), .B(G38), .ZN(new_n410_));
  NOR2_X1   g0096(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g0097(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g0098(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g0099(.A(G154), .ZN(new_n414_));
  AOI21_X1  g0100(.A(new_n377_), .B1(G18), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g0101(.A(new_n415_), .B(G2253), .ZN(new_n416_));
  INV_X1    g0102(.A(new_n416_), .ZN(new_n417_));
  OAI21_X1  g0103(.A(new_n383_), .B1(new_n371_), .B2(G155), .ZN(new_n418_));
  INV_X1    g0104(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g0105(.A1(new_n419_), .A2(G2247), .ZN(new_n420_));
  INV_X1    g0106(.A(G2247), .ZN(new_n421_));
  NAND2_X1  g0107(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g0108(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g0109(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g0110(.A(new_n383_), .B1(new_n371_), .B2(G153), .ZN(new_n425_));
  XNOR2_X1  g0111(.A(new_n425_), .B(G2256), .ZN(new_n426_));
  OAI21_X1  g0112(.A(new_n383_), .B1(new_n371_), .B2(G156), .ZN(new_n427_));
  XNOR2_X1  g0113(.A(new_n427_), .B(G2239), .ZN(new_n428_));
  NOR4_X1   g0114(.A1(new_n417_), .A2(new_n424_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n429_));
  OAI21_X1  g0115(.A(new_n383_), .B1(new_n371_), .B2(G157), .ZN(new_n430_));
  XNOR2_X1  g0116(.A(new_n430_), .B(G2236), .ZN(new_n431_));
  INV_X1    g0117(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g0118(.A1(G18), .A2(G159), .ZN(new_n433_));
  INV_X1    g0119(.A(G144), .ZN(new_n434_));
  OAI21_X1  g0120(.A(new_n433_), .B1(new_n434_), .B2(G18), .ZN(new_n435_));
  NAND2_X1  g0121(.A1(new_n435_), .A2(G2224), .ZN(new_n436_));
  INV_X1    g0122(.A(G2224), .ZN(new_n437_));
  OAI211_X1 g0123(.A(new_n433_), .B(new_n437_), .C1(G18), .C2(new_n434_), .ZN(new_n438_));
  NAND2_X1  g0124(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g0125(.A1(G18), .A2(G160), .ZN(new_n440_));
  INV_X1    g0126(.A(G138), .ZN(new_n441_));
  OAI21_X1  g0127(.A(new_n440_), .B1(new_n441_), .B2(G18), .ZN(new_n442_));
  NAND2_X1  g0128(.A1(new_n442_), .A2(G2218), .ZN(new_n443_));
  INV_X1    g0129(.A(G2218), .ZN(new_n444_));
  OAI211_X1 g0130(.A(new_n440_), .B(new_n444_), .C1(G18), .C2(new_n441_), .ZN(new_n445_));
  NAND2_X1  g0131(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g0132(.A1(new_n432_), .A2(new_n439_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g0133(.A1(new_n371_), .A2(G135), .ZN(new_n448_));
  INV_X1    g0134(.A(G158), .ZN(new_n449_));
  OAI21_X1  g0135(.A(new_n448_), .B1(new_n371_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g0136(.A1(new_n450_), .A2(G2230), .ZN(new_n451_));
  INV_X1    g0137(.A(G2230), .ZN(new_n452_));
  OAI211_X1 g0138(.A(new_n448_), .B(new_n452_), .C1(new_n371_), .C2(new_n449_), .ZN(new_n453_));
  NAND2_X1  g0139(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g0140(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g0141(.A1(new_n371_), .A2(G147), .ZN(new_n456_));
  NAND2_X1  g0142(.A1(G18), .A2(G151), .ZN(new_n457_));
  NAND2_X1  g0143(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g0144(.A(new_n458_), .B(G2211), .ZN(new_n459_));
  INV_X1    g0145(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g0146(.A1(new_n447_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  AND2_X1   g0147(.A1(new_n429_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g0148(.A1(new_n413_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g0149(.A1(new_n371_), .A2(G23), .ZN(new_n464_));
  INV_X1    g0150(.A(G236), .ZN(new_n465_));
  OAI21_X1  g0151(.A(new_n464_), .B1(new_n371_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g0152(.A1(new_n466_), .A2(G3717), .ZN(new_n467_));
  INV_X1    g0153(.A(G3717), .ZN(new_n468_));
  OAI211_X1 g0154(.A(new_n464_), .B(new_n468_), .C1(new_n371_), .C2(new_n465_), .ZN(new_n469_));
  NAND2_X1  g0155(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g0156(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g0157(.A(new_n372_), .ZN(new_n472_));
  NAND2_X1  g0158(.A1(new_n472_), .A2(new_n373_), .ZN(new_n473_));
  NOR2_X1   g0159(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g0160(.A1(G18), .A2(G237), .ZN(new_n475_));
  INV_X1    g0161(.A(G26), .ZN(new_n476_));
  OAI21_X1  g0162(.A(new_n475_), .B1(new_n476_), .B2(G18), .ZN(new_n477_));
  NAND2_X1  g0163(.A1(new_n477_), .A2(G3711), .ZN(new_n478_));
  INV_X1    g0164(.A(G3711), .ZN(new_n479_));
  OAI211_X1 g0165(.A(new_n475_), .B(new_n479_), .C1(G18), .C2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g0166(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g0167(.A1(G18), .A2(G238), .ZN(new_n482_));
  INV_X1    g0168(.A(G29), .ZN(new_n483_));
  OAI21_X1  g0169(.A(new_n482_), .B1(new_n483_), .B2(G18), .ZN(new_n484_));
  NAND2_X1  g0170(.A1(new_n484_), .A2(G3705), .ZN(new_n485_));
  INV_X1    g0171(.A(G3705), .ZN(new_n486_));
  OAI211_X1 g0172(.A(new_n482_), .B(new_n486_), .C1(G18), .C2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g0173(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g0174(.A1(new_n371_), .A2(G103), .ZN(new_n489_));
  INV_X1    g0175(.A(G235), .ZN(new_n490_));
  OAI21_X1  g0176(.A(new_n489_), .B1(new_n371_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g0177(.A(G3723), .ZN(new_n492_));
  XNOR2_X1  g0178(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g0179(.A(new_n493_), .ZN(new_n494_));
  NAND4_X1  g0180(.A1(new_n474_), .A2(new_n481_), .A3(new_n488_), .A4(new_n494_), .ZN(new_n495_));
  NAND2_X1  g0181(.A1(new_n491_), .A2(new_n492_), .ZN(new_n496_));
  NAND3_X1  g0182(.A1(new_n470_), .A2(new_n479_), .A3(new_n477_), .ZN(new_n497_));
  INV_X1    g0183(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g0184(.A1(new_n498_), .A2(new_n494_), .ZN(new_n499_));
  NAND2_X1  g0185(.A1(new_n371_), .A2(G29), .ZN(new_n500_));
  AOI21_X1  g0186(.A(G3705), .B1(new_n500_), .B2(new_n482_), .ZN(new_n501_));
  NAND4_X1  g0187(.A1(new_n494_), .A2(new_n470_), .A3(new_n481_), .A4(new_n501_), .ZN(new_n502_));
  NAND4_X1  g0188(.A1(new_n495_), .A2(new_n496_), .A3(new_n499_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g0189(.A1(new_n466_), .A2(new_n468_), .ZN(new_n504_));
  NOR2_X1   g0190(.A1(new_n493_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g0191(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g0192(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g0193(.A1(new_n371_), .A2(G124), .ZN(new_n508_));
  INV_X1    g0194(.A(G232), .ZN(new_n509_));
  OAI21_X1  g0195(.A(new_n508_), .B1(new_n371_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g0196(.A(new_n510_), .B(G3743), .ZN(new_n511_));
  INV_X1    g0197(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g0198(.A1(new_n371_), .A2(G127), .ZN(new_n513_));
  NAND2_X1  g0199(.A1(G18), .A2(G233), .ZN(new_n514_));
  NAND2_X1  g0200(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g0201(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g0202(.A(G3737), .ZN(new_n517_));
  NAND2_X1  g0203(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g0204(.A1(new_n515_), .A2(G3737), .ZN(new_n519_));
  NAND2_X1  g0205(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g0206(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g0207(.A1(new_n371_), .A2(G130), .ZN(new_n522_));
  INV_X1    g0208(.A(G234), .ZN(new_n523_));
  OAI21_X1  g0209(.A(new_n522_), .B1(new_n371_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g0210(.A(G3729), .ZN(new_n525_));
  XNOR2_X1  g0211(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g0212(.A1(new_n371_), .A2(G100), .ZN(new_n527_));
  INV_X1    g0213(.A(G231), .ZN(new_n528_));
  OAI21_X1  g0214(.A(new_n527_), .B1(new_n371_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g0215(.A(G3749), .ZN(new_n530_));
  XNOR2_X1  g0216(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR4_X1   g0217(.A1(new_n512_), .A2(new_n521_), .A3(new_n526_), .A4(new_n531_), .ZN(new_n532_));
  NAND2_X1  g0218(.A1(new_n507_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g0219(.A(new_n531_), .ZN(new_n534_));
  INV_X1    g0220(.A(new_n524_), .ZN(new_n535_));
  NOR2_X1   g0221(.A1(new_n535_), .A2(G3729), .ZN(new_n536_));
  INV_X1    g0222(.A(new_n536_), .ZN(new_n537_));
  NOR3_X1   g0223(.A1(new_n512_), .A2(new_n521_), .A3(new_n537_), .ZN(new_n538_));
  NOR2_X1   g0224(.A1(new_n516_), .A2(G3737), .ZN(new_n539_));
  NAND2_X1  g0225(.A1(new_n511_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g0226(.A(new_n540_), .ZN(new_n541_));
  OAI21_X1  g0227(.A(new_n534_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g0228(.A(G3743), .ZN(new_n543_));
  NAND2_X1  g0229(.A1(new_n510_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g0230(.A1(new_n531_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g0231(.A1(new_n529_), .A2(new_n530_), .ZN(new_n546_));
  NAND3_X1  g0232(.A1(new_n542_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g0233(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g0234(.A(new_n463_), .B1(new_n533_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g0235(.A1(new_n371_), .A2(G50), .ZN(new_n550_));
  INV_X1    g0236(.A(G220), .ZN(new_n551_));
  OAI21_X1  g0237(.A(new_n550_), .B1(new_n371_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g0238(.A(new_n552_), .B(G4432), .ZN(new_n553_));
  INV_X1    g0239(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g0240(.A1(new_n371_), .A2(G32), .ZN(new_n555_));
  NAND2_X1  g0241(.A1(G18), .A2(G221), .ZN(new_n556_));
  NAND2_X1  g0242(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g0243(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g0244(.A(G4427), .ZN(new_n559_));
  NAND2_X1  g0245(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g0246(.A1(new_n557_), .A2(G4427), .ZN(new_n561_));
  NAND2_X1  g0247(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g0248(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g0249(.A1(new_n371_), .A2(G66), .ZN(new_n564_));
  INV_X1    g0250(.A(G219), .ZN(new_n565_));
  OAI21_X1  g0251(.A(new_n564_), .B1(new_n371_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g0252(.A(G4437), .ZN(new_n567_));
  XNOR2_X1  g0253(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g0254(.A1(new_n371_), .A2(G35), .ZN(new_n569_));
  INV_X1    g0255(.A(G222), .ZN(new_n570_));
  OAI21_X1  g0256(.A(new_n569_), .B1(new_n371_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g0257(.A(G4420), .ZN(new_n572_));
  XNOR2_X1  g0258(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NOR4_X1   g0259(.A1(new_n554_), .A2(new_n563_), .A3(new_n568_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g0260(.A1(new_n371_), .A2(G47), .ZN(new_n575_));
  INV_X1    g0261(.A(G223), .ZN(new_n576_));
  OAI21_X1  g0262(.A(new_n575_), .B1(new_n371_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g0263(.A(new_n577_), .B(G4415), .ZN(new_n578_));
  NAND2_X1  g0264(.A1(new_n371_), .A2(G121), .ZN(new_n579_));
  INV_X1    g0265(.A(G224), .ZN(new_n580_));
  OAI21_X1  g0266(.A(new_n579_), .B1(new_n371_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g0267(.A1(new_n581_), .A2(G4410), .ZN(new_n582_));
  INV_X1    g0268(.A(G4410), .ZN(new_n583_));
  OAI211_X1 g0269(.A(new_n579_), .B(new_n583_), .C1(new_n371_), .C2(new_n580_), .ZN(new_n584_));
  NAND2_X1  g0270(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g0271(.A1(G18), .A2(G225), .ZN(new_n586_));
  INV_X1    g0272(.A(G94), .ZN(new_n587_));
  OAI21_X1  g0273(.A(new_n586_), .B1(new_n587_), .B2(G18), .ZN(new_n588_));
  NAND2_X1  g0274(.A1(new_n588_), .A2(G4405), .ZN(new_n589_));
  INV_X1    g0275(.A(G4405), .ZN(new_n590_));
  OAI211_X1 g0276(.A(new_n586_), .B(new_n590_), .C1(G18), .C2(new_n587_), .ZN(new_n591_));
  NAND2_X1  g0277(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g0278(.A1(G18), .A2(G226), .ZN(new_n593_));
  INV_X1    g0279(.A(G97), .ZN(new_n594_));
  OAI21_X1  g0280(.A(new_n593_), .B1(new_n594_), .B2(G18), .ZN(new_n595_));
  NAND2_X1  g0281(.A1(new_n595_), .A2(G4400), .ZN(new_n596_));
  INV_X1    g0282(.A(G4400), .ZN(new_n597_));
  OAI211_X1 g0283(.A(new_n593_), .B(new_n597_), .C1(G18), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g0284(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g0285(.A1(new_n578_), .A2(new_n585_), .A3(new_n592_), .A4(new_n599_), .ZN(new_n600_));
  NAND2_X1  g0286(.A1(new_n371_), .A2(G118), .ZN(new_n601_));
  NAND2_X1  g0287(.A1(G18), .A2(G217), .ZN(new_n602_));
  NAND2_X1  g0288(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g0289(.A(new_n603_), .B(G4394), .ZN(new_n604_));
  INV_X1    g0290(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g0291(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g0292(.A1(new_n574_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g0293(.A(new_n607_), .ZN(new_n608_));
  NOR3_X1   g0294(.A1(new_n463_), .A2(new_n375_), .A3(new_n607_), .ZN(new_n609_));
  NAND4_X1  g0295(.A1(new_n494_), .A2(new_n470_), .A3(new_n481_), .A4(new_n488_), .ZN(new_n610_));
  INV_X1    g0296(.A(new_n374_), .ZN(new_n611_));
  NOR2_X1   g0297(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g0298(.A1(new_n612_), .A2(new_n532_), .ZN(new_n613_));
  AOI22_X1  g0299(.A1(new_n549_), .A2(new_n608_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g0300(.A(new_n427_), .ZN(new_n615_));
  INV_X1    g0301(.A(G2239), .ZN(new_n616_));
  NAND2_X1  g0302(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g0303(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g0304(.A1(new_n416_), .A2(new_n423_), .A3(new_n618_), .ZN(new_n619_));
  NAND3_X1  g0305(.A1(new_n416_), .A2(new_n421_), .A3(new_n419_), .ZN(new_n620_));
  AOI21_X1  g0306(.A(new_n426_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g0307(.A(G2256), .ZN(new_n622_));
  INV_X1    g0308(.A(new_n425_), .ZN(new_n623_));
  AOI21_X1  g0309(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g0310(.A(G2253), .ZN(new_n625_));
  NAND2_X1  g0311(.A1(new_n415_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g0312(.A(new_n624_), .B1(new_n426_), .B2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g0313(.A(G2211), .B1(new_n456_), .B2(new_n457_), .ZN(new_n628_));
  INV_X1    g0314(.A(new_n628_), .ZN(new_n629_));
  NOR3_X1   g0315(.A1(new_n455_), .A2(new_n431_), .A3(new_n629_), .ZN(new_n630_));
  NAND3_X1  g0316(.A1(new_n630_), .A2(new_n439_), .A3(new_n446_), .ZN(new_n631_));
  OR2_X1    g0317(.A1(new_n430_), .A2(G2236), .ZN(new_n632_));
  NAND3_X1  g0318(.A1(new_n454_), .A2(new_n437_), .A3(new_n435_), .ZN(new_n633_));
  INV_X1    g0319(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g0320(.A1(new_n634_), .A2(new_n432_), .ZN(new_n635_));
  NAND2_X1  g0321(.A1(new_n371_), .A2(G138), .ZN(new_n636_));
  AOI21_X1  g0322(.A(G2218), .B1(new_n636_), .B2(new_n440_), .ZN(new_n637_));
  NAND4_X1  g0323(.A1(new_n432_), .A2(new_n454_), .A3(new_n439_), .A4(new_n637_), .ZN(new_n638_));
  NAND4_X1  g0324(.A1(new_n631_), .A2(new_n632_), .A3(new_n635_), .A4(new_n638_), .ZN(new_n639_));
  NAND2_X1  g0325(.A1(new_n450_), .A2(new_n452_), .ZN(new_n640_));
  NOR2_X1   g0326(.A1(new_n431_), .A2(new_n640_), .ZN(new_n641_));
  OR2_X1    g0327(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g0328(.A(new_n627_), .B1(new_n642_), .B2(new_n429_), .ZN(new_n643_));
  OR2_X1    g0329(.A1(new_n643_), .A2(new_n412_), .ZN(new_n644_));
  OAI21_X1  g0330(.A(G38), .B1(new_n407_), .B2(new_n409_), .ZN(new_n645_));
  INV_X1    g0331(.A(new_n645_), .ZN(new_n646_));
  OAI211_X1 g0332(.A(new_n383_), .B(new_n396_), .C1(new_n371_), .C2(G209), .ZN(new_n647_));
  NOR3_X1   g0333(.A1(new_n381_), .A2(new_n405_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g0334(.A1(new_n648_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n649_));
  NAND2_X1  g0335(.A1(new_n379_), .A2(new_n380_), .ZN(new_n650_));
  INV_X1    g0336(.A(G215), .ZN(new_n651_));
  NAND2_X1  g0337(.A1(new_n651_), .A2(G18), .ZN(new_n652_));
  NAND3_X1  g0338(.A1(new_n652_), .A2(new_n385_), .A3(new_n383_), .ZN(new_n653_));
  INV_X1    g0339(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g0340(.A1(new_n404_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g0341(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g0342(.A1(new_n656_), .A2(new_n382_), .ZN(new_n657_));
  INV_X1    g0343(.A(G216), .ZN(new_n658_));
  NAND2_X1  g0344(.A1(new_n658_), .A2(G18), .ZN(new_n659_));
  NAND3_X1  g0345(.A1(new_n659_), .A2(new_n390_), .A3(new_n383_), .ZN(new_n660_));
  INV_X1    g0346(.A(new_n660_), .ZN(new_n661_));
  NAND4_X1  g0347(.A1(new_n382_), .A2(new_n404_), .A3(new_n388_), .A4(new_n661_), .ZN(new_n662_));
  NAND4_X1  g0348(.A1(new_n649_), .A2(new_n650_), .A3(new_n657_), .A4(new_n662_), .ZN(new_n663_));
  NAND2_X1  g0349(.A1(new_n400_), .A2(new_n402_), .ZN(new_n664_));
  NOR2_X1   g0350(.A1(new_n381_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g0351(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g0352(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g0353(.A(new_n646_), .B1(new_n667_), .B2(new_n411_), .ZN(new_n668_));
  INV_X1    g0354(.A(new_n585_), .ZN(new_n669_));
  AOI21_X1  g0355(.A(G4394), .B1(new_n601_), .B2(new_n602_), .ZN(new_n670_));
  INV_X1    g0356(.A(new_n670_), .ZN(new_n671_));
  NOR2_X1   g0357(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g0358(.A1(new_n672_), .A2(new_n578_), .A3(new_n592_), .A4(new_n599_), .ZN(new_n673_));
  INV_X1    g0359(.A(G4415), .ZN(new_n674_));
  NAND2_X1  g0360(.A1(new_n577_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g0361(.A1(new_n585_), .A2(new_n590_), .A3(new_n588_), .ZN(new_n676_));
  INV_X1    g0362(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g0363(.A1(new_n677_), .A2(new_n578_), .ZN(new_n678_));
  NAND2_X1  g0364(.A1(new_n371_), .A2(G97), .ZN(new_n679_));
  AOI21_X1  g0365(.A(G4400), .B1(new_n679_), .B2(new_n593_), .ZN(new_n680_));
  NAND4_X1  g0366(.A1(new_n578_), .A2(new_n585_), .A3(new_n592_), .A4(new_n680_), .ZN(new_n681_));
  NAND4_X1  g0367(.A1(new_n673_), .A2(new_n675_), .A3(new_n678_), .A4(new_n681_), .ZN(new_n682_));
  INV_X1    g0368(.A(new_n578_), .ZN(new_n683_));
  NAND2_X1  g0369(.A1(new_n581_), .A2(new_n583_), .ZN(new_n684_));
  NOR2_X1   g0370(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OR2_X1    g0371(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g0372(.A1(new_n686_), .A2(new_n574_), .ZN(new_n687_));
  INV_X1    g0373(.A(G4432), .ZN(new_n688_));
  NAND2_X1  g0374(.A1(new_n552_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g0375(.A1(new_n568_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g0376(.A(new_n571_), .ZN(new_n691_));
  NOR2_X1   g0377(.A1(new_n691_), .A2(G4420), .ZN(new_n692_));
  NAND3_X1  g0378(.A1(new_n553_), .A2(new_n562_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g0379(.A1(new_n558_), .A2(G4427), .ZN(new_n694_));
  NAND2_X1  g0380(.A1(new_n553_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g0381(.A(new_n568_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  AOI211_X1 g0382(.A(new_n690_), .B(new_n696_), .C1(new_n567_), .C2(new_n566_), .ZN(new_n697_));
  NAND2_X1  g0383(.A1(new_n687_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g0384(.A1(new_n698_), .A2(new_n413_), .A3(new_n462_), .ZN(new_n699_));
  NAND4_X1  g0385(.A1(new_n614_), .A2(new_n644_), .A3(new_n668_), .A4(new_n699_), .ZN(G246));
  INV_X1    g0386(.A(G200), .ZN(new_n701_));
  OAI21_X1  g0387(.A(new_n527_), .B1(new_n371_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g0388(.A1(new_n371_), .A2(G56), .ZN(new_n703_));
  OAI21_X1  g0389(.A(new_n703_), .B1(new_n371_), .B2(G3749), .ZN(new_n704_));
  XOR2_X1   g0390(.A(new_n702_), .B(new_n704_), .Z(new_n705_));
  INV_X1    g0391(.A(G201), .ZN(new_n706_));
  OAI21_X1  g0392(.A(new_n508_), .B1(new_n371_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g0393(.A1(new_n371_), .A2(G55), .ZN(new_n708_));
  OAI21_X1  g0394(.A(new_n708_), .B1(new_n371_), .B2(G3743), .ZN(new_n709_));
  NAND3_X1  g0395(.A1(new_n705_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g0396(.A(G202), .ZN(new_n711_));
  OAI21_X1  g0397(.A(new_n513_), .B1(new_n371_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g0398(.A1(new_n371_), .A2(G54), .ZN(new_n713_));
  OAI21_X1  g0399(.A(new_n713_), .B1(new_n371_), .B2(G3737), .ZN(new_n714_));
  XOR2_X1   g0400(.A(new_n712_), .B(new_n714_), .Z(new_n715_));
  XOR2_X1   g0401(.A(new_n707_), .B(new_n709_), .Z(new_n716_));
  INV_X1    g0402(.A(new_n522_), .ZN(new_n717_));
  AOI21_X1  g0403(.A(new_n717_), .B1(G18), .B2(G203), .ZN(new_n718_));
  NOR2_X1   g0404(.A1(new_n371_), .A2(G3729), .ZN(new_n719_));
  AOI21_X1  g0405(.A(new_n719_), .B1(new_n371_), .B2(G53), .ZN(new_n720_));
  NOR2_X1   g0406(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g0407(.A1(new_n715_), .A2(new_n705_), .A3(new_n716_), .A4(new_n721_), .ZN(new_n722_));
  NAND4_X1  g0408(.A1(new_n705_), .A2(new_n716_), .A3(new_n712_), .A4(new_n714_), .ZN(new_n723_));
  NAND2_X1  g0409(.A1(new_n702_), .A2(new_n704_), .ZN(new_n724_));
  AND4_X1   g0410(.A1(new_n710_), .A2(new_n722_), .A3(new_n723_), .A4(new_n724_), .ZN(new_n725_));
  NAND2_X1  g0411(.A1(new_n371_), .A2(G41), .ZN(new_n726_));
  INV_X1    g0412(.A(G205), .ZN(new_n727_));
  OAI21_X1  g0413(.A(new_n464_), .B1(new_n371_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g0414(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g0415(.A1(new_n371_), .A2(G3717), .ZN(new_n730_));
  AOI21_X1  g0416(.A(new_n730_), .B1(new_n371_), .B2(G75), .ZN(new_n731_));
  XNOR2_X1  g0417(.A(new_n729_), .B(new_n731_), .ZN(new_n732_));
  INV_X1    g0418(.A(G70), .ZN(new_n733_));
  AOI211_X1 g0419(.A(new_n726_), .B(new_n732_), .C1(new_n371_), .C2(new_n733_), .ZN(new_n734_));
  INV_X1    g0420(.A(new_n500_), .ZN(new_n735_));
  AOI21_X1  g0421(.A(new_n735_), .B1(G18), .B2(G207), .ZN(new_n736_));
  NOR2_X1   g0422(.A1(new_n371_), .A2(G3705), .ZN(new_n737_));
  AOI21_X1  g0423(.A(new_n737_), .B1(new_n371_), .B2(G74), .ZN(new_n738_));
  XOR2_X1   g0424(.A(new_n736_), .B(new_n738_), .Z(new_n739_));
  NAND2_X1  g0425(.A1(new_n371_), .A2(G26), .ZN(new_n740_));
  INV_X1    g0426(.A(G206), .ZN(new_n741_));
  OAI21_X1  g0427(.A(new_n740_), .B1(new_n371_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g0428(.A1(new_n371_), .A2(G76), .ZN(new_n743_));
  OAI21_X1  g0429(.A(new_n743_), .B1(new_n371_), .B2(G3711), .ZN(new_n744_));
  XOR2_X1   g0430(.A(new_n742_), .B(new_n744_), .Z(new_n745_));
  NOR2_X1   g0431(.A1(new_n371_), .A2(G3723), .ZN(new_n746_));
  AOI21_X1  g0432(.A(new_n746_), .B1(new_n371_), .B2(G73), .ZN(new_n747_));
  INV_X1    g0433(.A(G204), .ZN(new_n748_));
  OAI21_X1  g0434(.A(new_n489_), .B1(new_n371_), .B2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g0435(.A(new_n747_), .B(new_n749_), .Z(new_n750_));
  INV_X1    g0436(.A(new_n750_), .ZN(new_n751_));
  NAND4_X1  g0437(.A1(new_n734_), .A2(new_n739_), .A3(new_n745_), .A4(new_n751_), .ZN(new_n752_));
  INV_X1    g0438(.A(new_n747_), .ZN(new_n753_));
  NAND2_X1  g0439(.A1(new_n753_), .A2(new_n749_), .ZN(new_n754_));
  INV_X1    g0440(.A(new_n732_), .ZN(new_n755_));
  NAND4_X1  g0441(.A1(new_n751_), .A2(new_n755_), .A3(new_n742_), .A4(new_n744_), .ZN(new_n756_));
  NOR3_X1   g0442(.A1(new_n732_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n757_));
  NAND3_X1  g0443(.A1(new_n757_), .A2(new_n745_), .A3(new_n751_), .ZN(new_n758_));
  NAND4_X1  g0444(.A1(new_n752_), .A2(new_n754_), .A3(new_n756_), .A4(new_n758_), .ZN(new_n759_));
  NOR3_X1   g0445(.A1(new_n750_), .A2(new_n729_), .A3(new_n731_), .ZN(new_n760_));
  NOR2_X1   g0446(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XOR2_X1   g0447(.A(new_n718_), .B(new_n720_), .Z(new_n762_));
  NAND4_X1  g0448(.A1(new_n762_), .A2(new_n715_), .A3(new_n705_), .A4(new_n716_), .ZN(new_n763_));
  OAI21_X1  g0449(.A(new_n725_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g0450(.A(new_n383_), .B1(new_n371_), .B2(G167), .ZN(new_n765_));
  INV_X1    g0451(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g0452(.A1(new_n371_), .A2(G112), .ZN(new_n767_));
  OAI21_X1  g0453(.A(new_n767_), .B1(new_n371_), .B2(G1480), .ZN(new_n768_));
  XNOR2_X1  g0454(.A(new_n766_), .B(new_n768_), .ZN(new_n769_));
  INV_X1    g0455(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g0456(.A(G166), .ZN(new_n771_));
  AOI21_X1  g0457(.A(new_n377_), .B1(G18), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g0458(.A1(new_n371_), .A2(G88), .ZN(new_n773_));
  OAI21_X1  g0459(.A(new_n773_), .B1(new_n371_), .B2(G1486), .ZN(new_n774_));
  XOR2_X1   g0460(.A(new_n772_), .B(new_n774_), .Z(new_n775_));
  NAND2_X1  g0461(.A1(new_n371_), .A2(G87), .ZN(new_n776_));
  OAI21_X1  g0462(.A(new_n776_), .B1(new_n371_), .B2(G106), .ZN(new_n777_));
  OAI21_X1  g0463(.A(new_n383_), .B1(new_n371_), .B2(G168), .ZN(new_n778_));
  XNOR2_X1  g0464(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  NAND3_X1  g0465(.A1(new_n770_), .A2(new_n775_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g0466(.A1(new_n371_), .A2(G111), .ZN(new_n781_));
  OAI21_X1  g0467(.A(new_n781_), .B1(new_n371_), .B2(G1469), .ZN(new_n782_));
  OAI21_X1  g0468(.A(new_n383_), .B1(new_n371_), .B2(G169), .ZN(new_n783_));
  XOR2_X1   g0469(.A(new_n782_), .B(new_n783_), .Z(new_n784_));
  NAND2_X1  g0470(.A1(new_n371_), .A2(G113), .ZN(new_n785_));
  OAI21_X1  g0471(.A(new_n785_), .B1(new_n371_), .B2(G1462), .ZN(new_n786_));
  XNOR2_X1  g0472(.A(new_n786_), .B(new_n383_), .ZN(new_n787_));
  NOR3_X1   g0473(.A1(new_n780_), .A2(new_n784_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g0474(.A(G4528), .ZN(new_n789_));
  NOR2_X1   g0475(.A1(new_n789_), .A2(G1455), .ZN(new_n790_));
  INV_X1    g0476(.A(G38), .ZN(new_n791_));
  XNOR2_X1  g0477(.A(new_n790_), .B(new_n791_), .ZN(new_n792_));
  NOR2_X1   g0478(.A1(new_n789_), .A2(G2204), .ZN(new_n793_));
  XNOR2_X1  g0479(.A(new_n793_), .B(new_n791_), .ZN(new_n794_));
  NOR2_X1   g0480(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  AND2_X1   g0481(.A1(new_n788_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g0482(.A(new_n448_), .ZN(new_n797_));
  AOI21_X1  g0483(.A(new_n797_), .B1(G18), .B2(G178), .ZN(new_n798_));
  NAND2_X1  g0484(.A1(new_n371_), .A2(G85), .ZN(new_n799_));
  OAI21_X1  g0485(.A(new_n799_), .B1(new_n371_), .B2(G2230), .ZN(new_n800_));
  INV_X1    g0486(.A(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g0487(.A(new_n798_), .B(new_n801_), .ZN(new_n802_));
  INV_X1    g0488(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g0489(.A1(new_n371_), .A2(G144), .ZN(new_n804_));
  INV_X1    g0490(.A(G179), .ZN(new_n805_));
  OAI21_X1  g0491(.A(new_n804_), .B1(new_n371_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g0492(.A1(new_n371_), .A2(G84), .ZN(new_n807_));
  OAI21_X1  g0493(.A(new_n807_), .B1(new_n371_), .B2(G2224), .ZN(new_n808_));
  XOR2_X1   g0494(.A(new_n806_), .B(new_n808_), .Z(new_n809_));
  INV_X1    g0495(.A(G171), .ZN(new_n810_));
  OAI21_X1  g0496(.A(new_n456_), .B1(new_n371_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g0497(.A1(new_n371_), .A2(G65), .ZN(new_n812_));
  OAI21_X1  g0498(.A(new_n812_), .B1(new_n371_), .B2(G2211), .ZN(new_n813_));
  XOR2_X1   g0499(.A(new_n811_), .B(new_n813_), .Z(new_n814_));
  OAI21_X1  g0500(.A(new_n383_), .B1(new_n371_), .B2(G177), .ZN(new_n815_));
  INV_X1    g0501(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g0502(.A1(new_n371_), .A2(G64), .ZN(new_n817_));
  OAI21_X1  g0503(.A(new_n817_), .B1(new_n371_), .B2(G2236), .ZN(new_n818_));
  XNOR2_X1  g0504(.A(new_n816_), .B(new_n818_), .ZN(new_n819_));
  INV_X1    g0505(.A(new_n819_), .ZN(new_n820_));
  NAND4_X1  g0506(.A1(new_n803_), .A2(new_n809_), .A3(new_n814_), .A4(new_n820_), .ZN(new_n821_));
  NAND2_X1  g0507(.A1(new_n371_), .A2(G110), .ZN(new_n822_));
  OAI21_X1  g0508(.A(new_n822_), .B1(new_n371_), .B2(G2256), .ZN(new_n823_));
  OAI21_X1  g0509(.A(new_n383_), .B1(new_n371_), .B2(G173), .ZN(new_n824_));
  XNOR2_X1  g0510(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  NAND2_X1  g0511(.A1(new_n371_), .A2(G86), .ZN(new_n826_));
  OAI21_X1  g0512(.A(new_n826_), .B1(new_n371_), .B2(G2247), .ZN(new_n827_));
  OAI21_X1  g0513(.A(new_n383_), .B1(new_n371_), .B2(G175), .ZN(new_n828_));
  XNOR2_X1  g0514(.A(new_n827_), .B(new_n828_), .ZN(new_n829_));
  NAND2_X1  g0515(.A1(new_n371_), .A2(G109), .ZN(new_n830_));
  OAI21_X1  g0516(.A(new_n830_), .B1(new_n371_), .B2(G2253), .ZN(new_n831_));
  OAI21_X1  g0517(.A(new_n383_), .B1(new_n371_), .B2(G174), .ZN(new_n832_));
  XNOR2_X1  g0518(.A(new_n831_), .B(new_n832_), .ZN(new_n833_));
  NAND2_X1  g0519(.A1(new_n371_), .A2(G63), .ZN(new_n834_));
  OAI21_X1  g0520(.A(new_n834_), .B1(new_n371_), .B2(G2239), .ZN(new_n835_));
  OAI21_X1  g0521(.A(new_n383_), .B1(new_n371_), .B2(G176), .ZN(new_n836_));
  XNOR2_X1  g0522(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  NAND4_X1  g0523(.A1(new_n825_), .A2(new_n829_), .A3(new_n833_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1    g0524(.A(new_n636_), .ZN(new_n839_));
  AOI21_X1  g0525(.A(new_n839_), .B1(G18), .B2(G180), .ZN(new_n840_));
  NAND2_X1  g0526(.A1(new_n371_), .A2(G83), .ZN(new_n841_));
  OAI21_X1  g0527(.A(new_n841_), .B1(new_n371_), .B2(G2218), .ZN(new_n842_));
  INV_X1    g0528(.A(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g0529(.A(new_n840_), .B(new_n843_), .ZN(new_n844_));
  NOR3_X1   g0530(.A1(new_n821_), .A2(new_n838_), .A3(new_n844_), .ZN(new_n845_));
  AND3_X1   g0531(.A1(new_n764_), .A2(new_n796_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g0532(.A1(new_n371_), .A2(G4410), .ZN(new_n847_));
  AOI21_X1  g0533(.A(new_n847_), .B1(new_n371_), .B2(G81), .ZN(new_n848_));
  INV_X1    g0534(.A(G194), .ZN(new_n849_));
  OAI21_X1  g0535(.A(new_n579_), .B1(new_n371_), .B2(new_n849_), .ZN(new_n850_));
  XOR2_X1   g0536(.A(new_n848_), .B(new_n850_), .Z(new_n851_));
  INV_X1    g0537(.A(new_n851_), .ZN(new_n852_));
  INV_X1    g0538(.A(G193), .ZN(new_n853_));
  OAI21_X1  g0539(.A(new_n575_), .B1(new_n371_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g0540(.A1(new_n371_), .A2(G80), .ZN(new_n855_));
  OAI21_X1  g0541(.A(new_n855_), .B1(new_n371_), .B2(G4415), .ZN(new_n856_));
  XOR2_X1   g0542(.A(new_n854_), .B(new_n856_), .Z(new_n857_));
  NAND2_X1  g0543(.A1(new_n371_), .A2(G94), .ZN(new_n858_));
  INV_X1    g0544(.A(G195), .ZN(new_n859_));
  OAI21_X1  g0545(.A(new_n858_), .B1(new_n371_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g0546(.A1(new_n371_), .A2(G59), .ZN(new_n861_));
  OAI21_X1  g0547(.A(new_n861_), .B1(new_n371_), .B2(G4405), .ZN(new_n862_));
  XOR2_X1   g0548(.A(new_n860_), .B(new_n862_), .Z(new_n863_));
  NOR2_X1   g0549(.A1(new_n371_), .A2(G4394), .ZN(new_n864_));
  AOI21_X1  g0550(.A(new_n864_), .B1(new_n371_), .B2(G77), .ZN(new_n865_));
  INV_X1    g0551(.A(G187), .ZN(new_n866_));
  OAI21_X1  g0552(.A(new_n601_), .B1(new_n371_), .B2(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g0553(.A(new_n865_), .B(new_n867_), .ZN(new_n868_));
  NAND4_X1  g0554(.A1(new_n852_), .A2(new_n857_), .A3(new_n863_), .A4(new_n868_), .ZN(new_n869_));
  INV_X1    g0555(.A(new_n679_), .ZN(new_n870_));
  AOI21_X1  g0556(.A(new_n870_), .B1(G18), .B2(G196), .ZN(new_n871_));
  NOR2_X1   g0557(.A1(new_n371_), .A2(G4400), .ZN(new_n872_));
  AOI21_X1  g0558(.A(new_n872_), .B1(new_n371_), .B2(G78), .ZN(new_n873_));
  XNOR2_X1  g0559(.A(new_n871_), .B(new_n873_), .ZN(new_n874_));
  NOR2_X1   g0560(.A1(new_n869_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g0561(.A(new_n569_), .ZN(new_n876_));
  AOI21_X1  g0562(.A(new_n876_), .B1(G18), .B2(G192), .ZN(new_n877_));
  NOR2_X1   g0563(.A1(new_n371_), .A2(G4420), .ZN(new_n878_));
  AOI21_X1  g0564(.A(new_n878_), .B1(new_n371_), .B2(G79), .ZN(new_n879_));
  XOR2_X1   g0565(.A(new_n877_), .B(new_n879_), .Z(new_n880_));
  INV_X1    g0566(.A(G189), .ZN(new_n881_));
  OAI21_X1  g0567(.A(new_n564_), .B1(new_n371_), .B2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g0568(.A1(new_n371_), .A2(G62), .ZN(new_n883_));
  OAI21_X1  g0569(.A(new_n883_), .B1(new_n371_), .B2(G4437), .ZN(new_n884_));
  XOR2_X1   g0570(.A(new_n882_), .B(new_n884_), .Z(new_n885_));
  INV_X1    g0571(.A(G191), .ZN(new_n886_));
  OAI21_X1  g0572(.A(new_n555_), .B1(new_n371_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g0573(.A1(new_n371_), .A2(G60), .ZN(new_n888_));
  OAI21_X1  g0574(.A(new_n888_), .B1(new_n371_), .B2(G4427), .ZN(new_n889_));
  XOR2_X1   g0575(.A(new_n887_), .B(new_n889_), .Z(new_n890_));
  INV_X1    g0576(.A(G190), .ZN(new_n891_));
  OAI21_X1  g0577(.A(new_n550_), .B1(new_n371_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g0578(.A1(new_n371_), .A2(G61), .ZN(new_n893_));
  OAI21_X1  g0579(.A(new_n893_), .B1(new_n371_), .B2(G4432), .ZN(new_n894_));
  XOR2_X1   g0580(.A(new_n892_), .B(new_n894_), .Z(new_n895_));
  NAND4_X1  g0581(.A1(new_n880_), .A2(new_n885_), .A3(new_n890_), .A4(new_n895_), .ZN(new_n896_));
  INV_X1    g0582(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g0583(.A1(new_n875_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g0584(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g0585(.A1(new_n750_), .A2(new_n732_), .ZN(new_n900_));
  NAND2_X1  g0586(.A1(new_n371_), .A2(new_n733_), .ZN(new_n901_));
  XNOR2_X1  g0587(.A(new_n901_), .B(new_n726_), .ZN(new_n902_));
  NAND4_X1  g0588(.A1(new_n900_), .A2(new_n739_), .A3(new_n902_), .A4(new_n745_), .ZN(new_n903_));
  NOR2_X1   g0589(.A1(new_n903_), .A2(new_n763_), .ZN(new_n904_));
  AND4_X1   g0590(.A1(G89), .A2(new_n899_), .A3(new_n796_), .A4(new_n845_), .ZN(new_n905_));
  AOI22_X1  g0591(.A1(new_n846_), .A2(new_n899_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  AND3_X1   g0592(.A1(new_n803_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n907_));
  INV_X1    g0593(.A(new_n844_), .ZN(new_n908_));
  NAND4_X1  g0594(.A1(new_n907_), .A2(new_n820_), .A3(new_n809_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g0595(.A1(new_n816_), .A2(new_n818_), .ZN(new_n910_));
  NAND4_X1  g0596(.A1(new_n803_), .A2(new_n820_), .A3(new_n806_), .A4(new_n808_), .ZN(new_n911_));
  NOR3_X1   g0597(.A1(new_n802_), .A2(new_n840_), .A3(new_n843_), .ZN(new_n912_));
  NAND3_X1  g0598(.A1(new_n912_), .A2(new_n820_), .A3(new_n809_), .ZN(new_n913_));
  NAND4_X1  g0599(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .A4(new_n913_), .ZN(new_n914_));
  NOR3_X1   g0600(.A1(new_n819_), .A2(new_n798_), .A3(new_n801_), .ZN(new_n915_));
  NOR2_X1   g0601(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g0602(.A1(new_n916_), .A2(new_n838_), .ZN(new_n917_));
  INV_X1    g0603(.A(new_n835_), .ZN(new_n918_));
  NOR2_X1   g0604(.A1(new_n918_), .A2(new_n836_), .ZN(new_n919_));
  NAND4_X1  g0605(.A1(new_n825_), .A2(new_n829_), .A3(new_n833_), .A4(new_n919_), .ZN(new_n920_));
  INV_X1    g0606(.A(new_n828_), .ZN(new_n921_));
  NAND4_X1  g0607(.A1(new_n825_), .A2(new_n833_), .A3(new_n921_), .A4(new_n827_), .ZN(new_n922_));
  INV_X1    g0608(.A(new_n832_), .ZN(new_n923_));
  NAND3_X1  g0609(.A1(new_n825_), .A2(new_n923_), .A3(new_n831_), .ZN(new_n924_));
  INV_X1    g0610(.A(new_n824_), .ZN(new_n925_));
  NAND2_X1  g0611(.A1(new_n925_), .A2(new_n823_), .ZN(new_n926_));
  NAND4_X1  g0612(.A1(new_n920_), .A2(new_n922_), .A3(new_n924_), .A4(new_n926_), .ZN(new_n927_));
  OAI21_X1  g0613(.A(new_n796_), .B1(new_n917_), .B2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g0614(.A(new_n791_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n929_));
  INV_X1    g0615(.A(new_n786_), .ZN(new_n930_));
  NOR3_X1   g0616(.A1(new_n769_), .A2(new_n377_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g0617(.A(new_n784_), .ZN(new_n932_));
  NAND4_X1  g0618(.A1(new_n931_), .A2(new_n932_), .A3(new_n779_), .A4(new_n775_), .ZN(new_n933_));
  INV_X1    g0619(.A(new_n782_), .ZN(new_n934_));
  NOR3_X1   g0620(.A1(new_n769_), .A2(new_n783_), .A3(new_n934_), .ZN(new_n935_));
  NAND3_X1  g0621(.A1(new_n935_), .A2(new_n779_), .A3(new_n775_), .ZN(new_n936_));
  AND2_X1   g0622(.A1(new_n933_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g0623(.A1(new_n775_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n938_));
  NAND2_X1  g0624(.A1(new_n772_), .A2(new_n774_), .ZN(new_n939_));
  INV_X1    g0625(.A(new_n778_), .ZN(new_n940_));
  NAND4_X1  g0626(.A1(new_n770_), .A2(new_n775_), .A3(new_n940_), .A4(new_n777_), .ZN(new_n941_));
  NAND4_X1  g0627(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .A4(new_n941_), .ZN(new_n942_));
  AOI21_X1  g0628(.A(new_n929_), .B1(new_n942_), .B2(new_n795_), .ZN(new_n943_));
  INV_X1    g0629(.A(new_n867_), .ZN(new_n944_));
  NOR3_X1   g0630(.A1(new_n851_), .A2(new_n944_), .A3(new_n865_), .ZN(new_n945_));
  INV_X1    g0631(.A(new_n874_), .ZN(new_n946_));
  NAND4_X1  g0632(.A1(new_n945_), .A2(new_n857_), .A3(new_n863_), .A4(new_n946_), .ZN(new_n947_));
  NOR3_X1   g0633(.A1(new_n851_), .A2(new_n871_), .A3(new_n873_), .ZN(new_n948_));
  NAND3_X1  g0634(.A1(new_n948_), .A2(new_n857_), .A3(new_n863_), .ZN(new_n949_));
  AND2_X1   g0635(.A1(new_n947_), .A2(new_n949_), .ZN(new_n950_));
  INV_X1    g0636(.A(new_n848_), .ZN(new_n951_));
  NAND3_X1  g0637(.A1(new_n857_), .A2(new_n850_), .A3(new_n951_), .ZN(new_n952_));
  NAND2_X1  g0638(.A1(new_n854_), .A2(new_n856_), .ZN(new_n953_));
  NAND4_X1  g0639(.A1(new_n852_), .A2(new_n857_), .A3(new_n860_), .A4(new_n862_), .ZN(new_n954_));
  NAND4_X1  g0640(.A1(new_n950_), .A2(new_n952_), .A3(new_n953_), .A4(new_n954_), .ZN(new_n955_));
  NAND2_X1  g0641(.A1(new_n955_), .A2(new_n897_), .ZN(new_n956_));
  NAND3_X1  g0642(.A1(new_n885_), .A2(new_n892_), .A3(new_n894_), .ZN(new_n957_));
  NOR2_X1   g0643(.A1(new_n877_), .A2(new_n879_), .ZN(new_n958_));
  NAND4_X1  g0644(.A1(new_n885_), .A2(new_n890_), .A3(new_n895_), .A4(new_n958_), .ZN(new_n959_));
  NAND4_X1  g0645(.A1(new_n885_), .A2(new_n895_), .A3(new_n887_), .A4(new_n889_), .ZN(new_n960_));
  NAND2_X1  g0646(.A1(new_n882_), .A2(new_n884_), .ZN(new_n961_));
  AND4_X1   g0647(.A1(new_n957_), .A2(new_n959_), .A3(new_n960_), .A4(new_n961_), .ZN(new_n962_));
  NAND2_X1  g0648(.A1(new_n956_), .A2(new_n962_), .ZN(new_n963_));
  NAND3_X1  g0649(.A1(new_n963_), .A2(new_n796_), .A3(new_n845_), .ZN(new_n964_));
  NAND4_X1  g0650(.A1(new_n906_), .A2(new_n928_), .A3(new_n943_), .A4(new_n964_), .ZN(G258));
  NAND4_X1  g0651(.A1(new_n906_), .A2(new_n928_), .A3(new_n943_), .A4(new_n964_), .ZN(G264));
  INV_X1    g0652(.A(new_n526_), .ZN(new_n967_));
  NAND4_X1  g0653(.A1(new_n967_), .A2(new_n534_), .A3(new_n511_), .A4(new_n520_), .ZN(new_n968_));
  OAI21_X1  g0654(.A(new_n548_), .B1(new_n506_), .B2(new_n968_), .ZN(new_n969_));
  INV_X1    g0655(.A(new_n969_), .ZN(new_n970_));
  INV_X1    g0656(.A(new_n591_), .ZN(new_n971_));
  AOI21_X1  g0657(.A(new_n590_), .B1(new_n858_), .B2(new_n586_), .ZN(new_n972_));
  NOR2_X1   g0658(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  NOR3_X1   g0659(.A1(new_n683_), .A2(new_n669_), .A3(new_n973_), .ZN(new_n974_));
  NAND3_X1  g0660(.A1(new_n974_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n975_));
  INV_X1    g0661(.A(new_n568_), .ZN(new_n976_));
  INV_X1    g0662(.A(new_n573_), .ZN(new_n977_));
  NAND4_X1  g0663(.A1(new_n976_), .A2(new_n977_), .A3(new_n562_), .A4(new_n553_), .ZN(new_n978_));
  NOR2_X1   g0664(.A1(new_n975_), .A2(new_n978_), .ZN(new_n979_));
  INV_X1    g0665(.A(new_n979_), .ZN(new_n980_));
  NAND4_X1  g0666(.A1(new_n382_), .A2(new_n397_), .A3(new_n404_), .A4(new_n388_), .ZN(new_n981_));
  INV_X1    g0667(.A(new_n393_), .ZN(new_n982_));
  NOR2_X1   g0668(.A1(new_n981_), .A2(new_n982_), .ZN(new_n983_));
  INV_X1    g0669(.A(new_n983_), .ZN(new_n984_));
  INV_X1    g0670(.A(new_n411_), .ZN(new_n985_));
  NOR2_X1   g0671(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  NOR4_X1   g0672(.A1(new_n417_), .A2(new_n424_), .A3(new_n426_), .A4(new_n428_), .ZN(new_n987_));
  NAND4_X1  g0673(.A1(new_n432_), .A2(new_n454_), .A3(new_n459_), .A4(new_n439_), .ZN(new_n988_));
  INV_X1    g0674(.A(new_n446_), .ZN(new_n989_));
  NOR2_X1   g0675(.A1(new_n988_), .A2(new_n989_), .ZN(new_n990_));
  AND2_X1   g0676(.A1(new_n987_), .A2(new_n990_), .ZN(new_n991_));
  NAND2_X1  g0677(.A1(new_n986_), .A2(new_n991_), .ZN(new_n992_));
  NOR3_X1   g0678(.A1(new_n970_), .A2(new_n980_), .A3(new_n992_), .ZN(new_n993_));
  NAND4_X1  g0679(.A1(new_n494_), .A2(new_n374_), .A3(new_n470_), .A4(new_n481_), .ZN(new_n994_));
  INV_X1    g0680(.A(new_n488_), .ZN(new_n995_));
  NOR2_X1   g0681(.A1(new_n994_), .A2(new_n995_), .ZN(new_n996_));
  INV_X1    g0682(.A(new_n996_), .ZN(new_n997_));
  NOR2_X1   g0683(.A1(new_n997_), .A2(new_n968_), .ZN(new_n998_));
  NOR3_X1   g0684(.A1(new_n992_), .A2(new_n375_), .A3(new_n980_), .ZN(new_n999_));
  AOI21_X1  g0685(.A(new_n993_), .B1(new_n998_), .B2(new_n999_), .ZN(new_n1000_));
  AND2_X1   g0686(.A1(new_n642_), .A2(new_n987_), .ZN(new_n1001_));
  OAI21_X1  g0687(.A(new_n986_), .B1(new_n1001_), .B2(new_n627_), .ZN(new_n1002_));
  INV_X1    g0688(.A(new_n978_), .ZN(new_n1003_));
  NAND2_X1  g0689(.A1(new_n686_), .A2(new_n1003_), .ZN(new_n1004_));
  NAND2_X1  g0690(.A1(new_n1004_), .A2(new_n697_), .ZN(new_n1005_));
  NAND3_X1  g0691(.A1(new_n1005_), .A2(new_n986_), .A3(new_n991_), .ZN(new_n1006_));
  NAND4_X1  g0692(.A1(new_n1000_), .A2(new_n668_), .A3(new_n1002_), .A4(new_n1006_), .ZN(G270));
  NAND3_X1  g0693(.A1(new_n470_), .A2(new_n481_), .A3(new_n501_), .ZN(new_n1008_));
  AOI21_X1  g0694(.A(new_n372_), .B1(new_n371_), .B2(G3701), .ZN(new_n1009_));
  NAND4_X1  g0695(.A1(new_n470_), .A2(new_n481_), .A3(new_n488_), .A4(new_n1009_), .ZN(new_n1010_));
  NAND4_X1  g0696(.A1(new_n470_), .A2(G4526), .A3(new_n481_), .A4(new_n488_), .ZN(new_n1011_));
  OAI211_X1 g0697(.A(new_n1008_), .B(new_n1010_), .C1(new_n1011_), .C2(new_n611_), .ZN(new_n1012_));
  INV_X1    g0698(.A(new_n1012_), .ZN(new_n1013_));
  NAND3_X1  g0699(.A1(new_n1013_), .A2(new_n504_), .A3(new_n497_), .ZN(new_n1014_));
  XNOR2_X1  g0700(.A(new_n1014_), .B(new_n493_), .ZN(G388));
  AOI21_X1  g0701(.A(new_n473_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n1016_));
  NAND2_X1  g0702(.A1(new_n1016_), .A2(new_n481_), .ZN(new_n1017_));
  NAND4_X1  g0703(.A1(new_n374_), .A2(new_n481_), .A3(new_n488_), .A4(G4526), .ZN(new_n1018_));
  NAND2_X1  g0704(.A1(new_n477_), .A2(new_n479_), .ZN(new_n1019_));
  INV_X1    g0705(.A(new_n480_), .ZN(new_n1020_));
  AOI21_X1  g0706(.A(new_n479_), .B1(new_n740_), .B2(new_n475_), .ZN(new_n1021_));
  OAI21_X1  g0707(.A(new_n501_), .B1(new_n1020_), .B2(new_n1021_), .ZN(new_n1022_));
  NAND4_X1  g0708(.A1(new_n1017_), .A2(new_n1018_), .A3(new_n1019_), .A4(new_n1022_), .ZN(new_n1023_));
  XNOR2_X1  g0709(.A(new_n1023_), .B(new_n471_), .ZN(G391));
  NAND3_X1  g0710(.A1(new_n374_), .A2(new_n488_), .A3(G4526), .ZN(new_n1025_));
  INV_X1    g0711(.A(new_n501_), .ZN(new_n1026_));
  INV_X1    g0712(.A(new_n487_), .ZN(new_n1027_));
  AOI21_X1  g0713(.A(new_n486_), .B1(new_n500_), .B2(new_n482_), .ZN(new_n1028_));
  OAI21_X1  g0714(.A(new_n1009_), .B1(new_n1027_), .B2(new_n1028_), .ZN(new_n1029_));
  NAND3_X1  g0715(.A1(new_n1025_), .A2(new_n1026_), .A3(new_n1029_), .ZN(new_n1030_));
  NOR2_X1   g0716(.A1(new_n1020_), .A2(new_n1021_), .ZN(new_n1031_));
  XNOR2_X1  g0717(.A(new_n1030_), .B(new_n1031_), .ZN(G394));
  AOI21_X1  g0718(.A(new_n1009_), .B1(new_n374_), .B2(G4526), .ZN(new_n1033_));
  XNOR2_X1  g0719(.A(new_n1033_), .B(new_n488_), .ZN(G397));
  AOI21_X1  g0720(.A(new_n507_), .B1(G4526), .B2(new_n612_), .ZN(new_n1035_));
  INV_X1    g0721(.A(new_n538_), .ZN(new_n1036_));
  NAND3_X1  g0722(.A1(new_n1036_), .A2(new_n544_), .A3(new_n540_), .ZN(new_n1037_));
  XNOR2_X1  g0723(.A(new_n1037_), .B(new_n531_), .ZN(new_n1038_));
  NAND2_X1  g0724(.A1(new_n1035_), .A2(new_n1038_), .ZN(new_n1039_));
  OAI211_X1 g0725(.A(new_n511_), .B(new_n520_), .C1(new_n525_), .C2(new_n524_), .ZN(new_n1040_));
  NAND3_X1  g0726(.A1(new_n1040_), .A2(new_n544_), .A3(new_n540_), .ZN(new_n1041_));
  XNOR2_X1  g0727(.A(new_n1041_), .B(new_n534_), .ZN(new_n1042_));
  OAI21_X1  g0728(.A(new_n1039_), .B1(new_n1035_), .B2(new_n1042_), .ZN(G376));
  NAND2_X1  g0729(.A1(new_n520_), .A2(new_n536_), .ZN(new_n1044_));
  INV_X1    g0730(.A(new_n539_), .ZN(new_n1045_));
  NAND2_X1  g0731(.A1(new_n1044_), .A2(new_n1045_), .ZN(new_n1046_));
  XNOR2_X1  g0732(.A(new_n1046_), .B(new_n512_), .ZN(new_n1047_));
  NAND2_X1  g0733(.A1(new_n1035_), .A2(new_n1047_), .ZN(new_n1048_));
  OAI211_X1 g0734(.A(new_n1044_), .B(new_n1045_), .C1(new_n521_), .C2(new_n526_), .ZN(new_n1049_));
  XNOR2_X1  g0735(.A(new_n1049_), .B(new_n511_), .ZN(new_n1050_));
  OAI21_X1  g0736(.A(new_n1048_), .B1(new_n1035_), .B2(new_n1050_), .ZN(G379));
  XNOR2_X1  g0737(.A(new_n537_), .B(new_n520_), .ZN(new_n1052_));
  NAND2_X1  g0738(.A1(new_n1035_), .A2(new_n1052_), .ZN(new_n1053_));
  NAND2_X1  g0739(.A1(new_n535_), .A2(G3729), .ZN(new_n1054_));
  XNOR2_X1  g0740(.A(new_n520_), .B(new_n1054_), .ZN(new_n1055_));
  OAI21_X1  g0741(.A(new_n1053_), .B1(new_n1035_), .B2(new_n1055_), .ZN(G382));
  XNOR2_X1  g0742(.A(new_n1035_), .B(new_n967_), .ZN(G385));
  XOR2_X1   g0743(.A(new_n450_), .B(new_n430_), .Z(new_n1058_));
  INV_X1    g0744(.A(new_n1058_), .ZN(new_n1059_));
  NAND2_X1  g0745(.A1(new_n371_), .A2(G141), .ZN(new_n1060_));
  INV_X1    g0746(.A(G161), .ZN(new_n1061_));
  OAI21_X1  g0747(.A(new_n1060_), .B1(new_n371_), .B2(new_n1061_), .ZN(new_n1062_));
  XNOR2_X1  g0748(.A(new_n1062_), .B(new_n458_), .ZN(new_n1063_));
  XNOR2_X1  g0749(.A(new_n435_), .B(new_n442_), .ZN(new_n1064_));
  NAND3_X1  g0750(.A1(new_n1059_), .A2(new_n1063_), .A3(new_n1064_), .ZN(new_n1065_));
  INV_X1    g0751(.A(new_n1064_), .ZN(new_n1066_));
  INV_X1    g0752(.A(new_n1063_), .ZN(new_n1067_));
  NAND3_X1  g0753(.A1(new_n1059_), .A2(new_n1066_), .A3(new_n1067_), .ZN(new_n1068_));
  NAND3_X1  g0754(.A1(new_n1067_), .A2(new_n1058_), .A3(new_n1064_), .ZN(new_n1069_));
  NAND3_X1  g0755(.A1(new_n1058_), .A2(new_n1066_), .A3(new_n1063_), .ZN(new_n1070_));
  NAND4_X1  g0756(.A1(new_n1065_), .A2(new_n1068_), .A3(new_n1069_), .A4(new_n1070_), .ZN(new_n1071_));
  XNOR2_X1  g0757(.A(new_n415_), .B(new_n425_), .ZN(new_n1072_));
  XOR2_X1   g0758(.A(new_n418_), .B(new_n427_), .Z(new_n1073_));
  XNOR2_X1  g0759(.A(new_n1072_), .B(new_n1073_), .ZN(new_n1074_));
  XNOR2_X1  g0760(.A(new_n1071_), .B(new_n1074_), .ZN(new_n1075_));
  OR2_X1    g0761(.A1(new_n379_), .A2(new_n399_), .ZN(new_n1076_));
  NAND2_X1  g0762(.A1(new_n379_), .A2(new_n399_), .ZN(new_n1077_));
  NAND2_X1  g0763(.A1(new_n1076_), .A2(new_n1077_), .ZN(new_n1078_));
  INV_X1    g0764(.A(new_n1078_), .ZN(new_n1079_));
  XNOR2_X1  g0765(.A(new_n384_), .B(new_n389_), .ZN(new_n1080_));
  NOR3_X1   g0766(.A1(new_n377_), .A2(new_n371_), .A3(G209), .ZN(new_n1081_));
  INV_X1    g0767(.A(new_n1081_), .ZN(new_n1082_));
  NAND3_X1  g0768(.A1(new_n1079_), .A2(new_n1080_), .A3(new_n1082_), .ZN(new_n1083_));
  INV_X1    g0769(.A(new_n1080_), .ZN(new_n1084_));
  NAND3_X1  g0770(.A1(new_n1079_), .A2(new_n1084_), .A3(new_n1081_), .ZN(new_n1085_));
  NAND3_X1  g0771(.A1(new_n1078_), .A2(new_n1080_), .A3(new_n1081_), .ZN(new_n1086_));
  NAND3_X1  g0772(.A1(new_n1078_), .A2(new_n1084_), .A3(new_n1082_), .ZN(new_n1087_));
  NAND4_X1  g0773(.A1(new_n1083_), .A2(new_n1085_), .A3(new_n1086_), .A4(new_n1087_), .ZN(new_n1088_));
  OAI21_X1  g0774(.A(new_n383_), .B1(new_n371_), .B2(G212), .ZN(new_n1089_));
  OAI21_X1  g0775(.A(new_n383_), .B1(new_n371_), .B2(G211), .ZN(new_n1090_));
  XNOR2_X1  g0776(.A(new_n1089_), .B(new_n1090_), .ZN(new_n1091_));
  XNOR2_X1  g0777(.A(new_n1088_), .B(new_n1091_), .ZN(new_n1092_));
  XNOR2_X1  g0778(.A(new_n466_), .B(new_n491_), .ZN(new_n1093_));
  INV_X1    g0779(.A(new_n1093_), .ZN(new_n1094_));
  NAND2_X1  g0780(.A1(new_n371_), .A2(G41), .ZN(new_n1095_));
  INV_X1    g0781(.A(G229), .ZN(new_n1096_));
  OAI21_X1  g0782(.A(new_n1095_), .B1(new_n371_), .B2(new_n1096_), .ZN(new_n1097_));
  NAND2_X1  g0783(.A1(new_n371_), .A2(G44), .ZN(new_n1098_));
  INV_X1    g0784(.A(G239), .ZN(new_n1099_));
  OAI21_X1  g0785(.A(new_n1098_), .B1(new_n371_), .B2(new_n1099_), .ZN(new_n1100_));
  XNOR2_X1  g0786(.A(new_n1097_), .B(new_n1100_), .ZN(new_n1101_));
  INV_X1    g0787(.A(new_n1101_), .ZN(new_n1102_));
  XNOR2_X1  g0788(.A(new_n477_), .B(new_n484_), .ZN(new_n1103_));
  INV_X1    g0789(.A(new_n1103_), .ZN(new_n1104_));
  NAND3_X1  g0790(.A1(new_n1094_), .A2(new_n1102_), .A3(new_n1104_), .ZN(new_n1105_));
  NAND3_X1  g0791(.A1(new_n1102_), .A2(new_n1103_), .A3(new_n1093_), .ZN(new_n1106_));
  NAND3_X1  g0792(.A1(new_n1094_), .A2(new_n1103_), .A3(new_n1101_), .ZN(new_n1107_));
  NAND3_X1  g0793(.A1(new_n1104_), .A2(new_n1093_), .A3(new_n1101_), .ZN(new_n1108_));
  NAND4_X1  g0794(.A1(new_n1105_), .A2(new_n1106_), .A3(new_n1107_), .A4(new_n1108_), .ZN(new_n1109_));
  XNOR2_X1  g0795(.A(new_n510_), .B(new_n529_), .ZN(new_n1110_));
  XNOR2_X1  g0796(.A(new_n524_), .B(new_n515_), .ZN(new_n1111_));
  XNOR2_X1  g0797(.A(new_n1110_), .B(new_n1111_), .ZN(new_n1112_));
  XNOR2_X1  g0798(.A(new_n1109_), .B(new_n1112_), .ZN(new_n1113_));
  XNOR2_X1  g0799(.A(new_n577_), .B(new_n581_), .ZN(new_n1114_));
  INV_X1    g0800(.A(new_n1114_), .ZN(new_n1115_));
  XNOR2_X1  g0801(.A(new_n588_), .B(new_n595_), .ZN(new_n1116_));
  NAND2_X1  g0802(.A1(new_n371_), .A2(G115), .ZN(new_n1117_));
  INV_X1    g0803(.A(G227), .ZN(new_n1118_));
  OAI21_X1  g0804(.A(new_n1117_), .B1(new_n371_), .B2(new_n1118_), .ZN(new_n1119_));
  XNOR2_X1  g0805(.A(new_n1119_), .B(new_n603_), .ZN(new_n1120_));
  NAND3_X1  g0806(.A1(new_n1115_), .A2(new_n1116_), .A3(new_n1120_), .ZN(new_n1121_));
  INV_X1    g0807(.A(new_n1120_), .ZN(new_n1122_));
  INV_X1    g0808(.A(new_n1116_), .ZN(new_n1123_));
  NAND3_X1  g0809(.A1(new_n1115_), .A2(new_n1122_), .A3(new_n1123_), .ZN(new_n1124_));
  NAND3_X1  g0810(.A1(new_n1122_), .A2(new_n1116_), .A3(new_n1114_), .ZN(new_n1125_));
  NAND3_X1  g0811(.A1(new_n1123_), .A2(new_n1114_), .A3(new_n1120_), .ZN(new_n1126_));
  NAND4_X1  g0812(.A1(new_n1121_), .A2(new_n1124_), .A3(new_n1125_), .A4(new_n1126_), .ZN(new_n1127_));
  XNOR2_X1  g0813(.A(new_n566_), .B(new_n552_), .ZN(new_n1128_));
  XNOR2_X1  g0814(.A(new_n571_), .B(new_n557_), .ZN(new_n1129_));
  XNOR2_X1  g0815(.A(new_n1128_), .B(new_n1129_), .ZN(new_n1130_));
  XNOR2_X1  g0816(.A(new_n1127_), .B(new_n1130_), .ZN(new_n1131_));
  NAND4_X1  g0817(.A1(new_n1075_), .A2(new_n1092_), .A3(new_n1113_), .A4(new_n1131_), .ZN(G412));
  XOR2_X1   g0818(.A(new_n738_), .B(new_n744_), .Z(new_n1133_));
  INV_X1    g0819(.A(new_n1133_), .ZN(new_n1134_));
  NOR2_X1   g0820(.A1(new_n371_), .A2(G3698), .ZN(new_n1135_));
  AOI21_X1  g0821(.A(new_n1135_), .B1(new_n371_), .B2(G69), .ZN(new_n1136_));
  NAND2_X1  g0822(.A1(new_n371_), .A2(G70), .ZN(new_n1137_));
  OAI21_X1  g0823(.A(new_n1137_), .B1(new_n371_), .B2(G3701), .ZN(new_n1138_));
  XOR2_X1   g0824(.A(new_n1136_), .B(new_n1138_), .Z(new_n1139_));
  INV_X1    g0825(.A(new_n1139_), .ZN(new_n1140_));
  XNOR2_X1  g0826(.A(new_n747_), .B(new_n731_), .ZN(new_n1141_));
  INV_X1    g0827(.A(new_n1141_), .ZN(new_n1142_));
  NAND3_X1  g0828(.A1(new_n1134_), .A2(new_n1140_), .A3(new_n1142_), .ZN(new_n1143_));
  NAND3_X1  g0829(.A1(new_n1140_), .A2(new_n1133_), .A3(new_n1141_), .ZN(new_n1144_));
  NAND3_X1  g0830(.A1(new_n1134_), .A2(new_n1141_), .A3(new_n1139_), .ZN(new_n1145_));
  NAND3_X1  g0831(.A1(new_n1142_), .A2(new_n1133_), .A3(new_n1139_), .ZN(new_n1146_));
  NAND4_X1  g0832(.A1(new_n1143_), .A2(new_n1144_), .A3(new_n1145_), .A4(new_n1146_), .ZN(new_n1147_));
  XOR2_X1   g0833(.A(new_n704_), .B(new_n709_), .Z(new_n1148_));
  XNOR2_X1  g0834(.A(new_n720_), .B(new_n714_), .ZN(new_n1149_));
  XNOR2_X1  g0835(.A(new_n1148_), .B(new_n1149_), .ZN(new_n1150_));
  XNOR2_X1  g0836(.A(new_n1147_), .B(new_n1150_), .ZN(new_n1151_));
  XOR2_X1   g0837(.A(new_n873_), .B(new_n862_), .Z(new_n1152_));
  INV_X1    g0838(.A(new_n1152_), .ZN(new_n1153_));
  XOR2_X1   g0839(.A(new_n848_), .B(new_n856_), .Z(new_n1154_));
  INV_X1    g0840(.A(new_n1154_), .ZN(new_n1155_));
  NOR2_X1   g0841(.A1(new_n371_), .A2(G4393), .ZN(new_n1156_));
  AOI21_X1  g0842(.A(new_n1156_), .B1(new_n371_), .B2(G58), .ZN(new_n1157_));
  XNOR2_X1  g0843(.A(new_n865_), .B(new_n1157_), .ZN(new_n1158_));
  INV_X1    g0844(.A(new_n1158_), .ZN(new_n1159_));
  NAND3_X1  g0845(.A1(new_n1153_), .A2(new_n1155_), .A3(new_n1159_), .ZN(new_n1160_));
  NAND3_X1  g0846(.A1(new_n1155_), .A2(new_n1158_), .A3(new_n1152_), .ZN(new_n1161_));
  NAND3_X1  g0847(.A1(new_n1153_), .A2(new_n1158_), .A3(new_n1154_), .ZN(new_n1162_));
  NAND3_X1  g0848(.A1(new_n1159_), .A2(new_n1152_), .A3(new_n1154_), .ZN(new_n1163_));
  NAND4_X1  g0849(.A1(new_n1160_), .A2(new_n1161_), .A3(new_n1162_), .A4(new_n1163_), .ZN(new_n1164_));
  XOR2_X1   g0850(.A(new_n884_), .B(new_n894_), .Z(new_n1165_));
  XNOR2_X1  g0851(.A(new_n879_), .B(new_n889_), .ZN(new_n1166_));
  XNOR2_X1  g0852(.A(new_n1165_), .B(new_n1166_), .ZN(new_n1167_));
  XNOR2_X1  g0853(.A(new_n1164_), .B(new_n1167_), .ZN(new_n1168_));
  NOR2_X1   g0854(.A1(new_n371_), .A2(G2208), .ZN(new_n1169_));
  AOI21_X1  g0855(.A(new_n1169_), .B1(new_n371_), .B2(G82), .ZN(new_n1170_));
  XOR2_X1   g0856(.A(new_n1170_), .B(new_n813_), .Z(new_n1171_));
  INV_X1    g0857(.A(new_n1171_), .ZN(new_n1172_));
  XNOR2_X1  g0858(.A(new_n808_), .B(new_n842_), .ZN(new_n1173_));
  XNOR2_X1  g0859(.A(new_n818_), .B(new_n800_), .ZN(new_n1174_));
  NAND3_X1  g0860(.A1(new_n1172_), .A2(new_n1173_), .A3(new_n1174_), .ZN(new_n1175_));
  INV_X1    g0861(.A(new_n1173_), .ZN(new_n1176_));
  INV_X1    g0862(.A(new_n1174_), .ZN(new_n1177_));
  NAND3_X1  g0863(.A1(new_n1172_), .A2(new_n1176_), .A3(new_n1177_), .ZN(new_n1178_));
  NAND3_X1  g0864(.A1(new_n1171_), .A2(new_n1173_), .A3(new_n1177_), .ZN(new_n1179_));
  NAND3_X1  g0865(.A1(new_n1171_), .A2(new_n1176_), .A3(new_n1174_), .ZN(new_n1180_));
  NAND4_X1  g0866(.A1(new_n1175_), .A2(new_n1178_), .A3(new_n1179_), .A4(new_n1180_), .ZN(new_n1181_));
  XNOR2_X1  g0867(.A(new_n827_), .B(new_n835_), .ZN(new_n1182_));
  XNOR2_X1  g0868(.A(new_n823_), .B(new_n831_), .ZN(new_n1183_));
  XNOR2_X1  g0869(.A(new_n1182_), .B(new_n1183_), .ZN(new_n1184_));
  XNOR2_X1  g0870(.A(new_n1181_), .B(new_n1184_), .ZN(new_n1185_));
  NOR2_X1   g0871(.A1(new_n371_), .A2(G1459), .ZN(new_n1186_));
  AOI21_X1  g0872(.A(new_n1186_), .B1(new_n371_), .B2(G114), .ZN(new_n1187_));
  XNOR2_X1  g0873(.A(new_n930_), .B(new_n1187_), .ZN(new_n1188_));
  INV_X1    g0874(.A(new_n1188_), .ZN(new_n1189_));
  XNOR2_X1  g0875(.A(new_n782_), .B(new_n777_), .ZN(new_n1190_));
  XNOR2_X1  g0876(.A(new_n774_), .B(new_n768_), .ZN(new_n1191_));
  NAND3_X1  g0877(.A1(new_n1189_), .A2(new_n1190_), .A3(new_n1191_), .ZN(new_n1192_));
  INV_X1    g0878(.A(new_n1190_), .ZN(new_n1193_));
  INV_X1    g0879(.A(new_n1191_), .ZN(new_n1194_));
  NAND3_X1  g0880(.A1(new_n1189_), .A2(new_n1193_), .A3(new_n1194_), .ZN(new_n1195_));
  NAND3_X1  g0881(.A1(new_n1194_), .A2(new_n1188_), .A3(new_n1190_), .ZN(new_n1196_));
  NAND3_X1  g0882(.A1(new_n1193_), .A2(new_n1188_), .A3(new_n1191_), .ZN(new_n1197_));
  NAND4_X1  g0883(.A1(new_n1192_), .A2(new_n1195_), .A3(new_n1196_), .A4(new_n1197_), .ZN(new_n1198_));
  NAND2_X1  g0884(.A1(new_n371_), .A2(G1455), .ZN(new_n1199_));
  OAI21_X1  g0885(.A(new_n1199_), .B1(new_n371_), .B2(G1492), .ZN(new_n1200_));
  NAND2_X1  g0886(.A1(new_n371_), .A2(G2204), .ZN(new_n1201_));
  OAI21_X1  g0887(.A(new_n1201_), .B1(new_n371_), .B2(G1496), .ZN(new_n1202_));
  XNOR2_X1  g0888(.A(new_n1200_), .B(new_n1202_), .ZN(new_n1203_));
  XNOR2_X1  g0889(.A(new_n1198_), .B(new_n1203_), .ZN(new_n1204_));
  NAND4_X1  g0890(.A1(new_n1151_), .A2(new_n1168_), .A3(new_n1185_), .A4(new_n1204_), .ZN(G414));
  XOR2_X1   g0891(.A(new_n840_), .B(new_n806_), .Z(new_n1206_));
  INV_X1    g0892(.A(new_n1206_), .ZN(new_n1207_));
  XNOR2_X1  g0893(.A(new_n798_), .B(new_n815_), .ZN(new_n1208_));
  INV_X1    g0894(.A(G181), .ZN(new_n1209_));
  OAI21_X1  g0895(.A(new_n1060_), .B1(new_n371_), .B2(new_n1209_), .ZN(new_n1210_));
  XNOR2_X1  g0896(.A(new_n811_), .B(new_n1210_), .ZN(new_n1211_));
  NAND3_X1  g0897(.A1(new_n1207_), .A2(new_n1208_), .A3(new_n1211_), .ZN(new_n1212_));
  INV_X1    g0898(.A(new_n1211_), .ZN(new_n1213_));
  INV_X1    g0899(.A(new_n1208_), .ZN(new_n1214_));
  NAND3_X1  g0900(.A1(new_n1207_), .A2(new_n1213_), .A3(new_n1214_), .ZN(new_n1215_));
  NAND3_X1  g0901(.A1(new_n1206_), .A2(new_n1208_), .A3(new_n1213_), .ZN(new_n1216_));
  NAND3_X1  g0902(.A1(new_n1214_), .A2(new_n1206_), .A3(new_n1211_), .ZN(new_n1217_));
  NAND4_X1  g0903(.A1(new_n1212_), .A2(new_n1215_), .A3(new_n1216_), .A4(new_n1217_), .ZN(new_n1218_));
  XNOR2_X1  g0904(.A(new_n828_), .B(new_n836_), .ZN(new_n1219_));
  XNOR2_X1  g0905(.A(new_n824_), .B(new_n832_), .ZN(new_n1220_));
  XNOR2_X1  g0906(.A(new_n1219_), .B(new_n1220_), .ZN(new_n1221_));
  XNOR2_X1  g0907(.A(new_n1218_), .B(new_n1221_), .ZN(new_n1222_));
  XOR2_X1   g0908(.A(new_n736_), .B(new_n742_), .Z(new_n1223_));
  INV_X1    g0909(.A(new_n1223_), .ZN(new_n1224_));
  XNOR2_X1  g0910(.A(new_n749_), .B(new_n728_), .ZN(new_n1225_));
  INV_X1    g0911(.A(G198), .ZN(new_n1226_));
  OAI21_X1  g0912(.A(new_n1095_), .B1(new_n371_), .B2(new_n1226_), .ZN(new_n1227_));
  INV_X1    g0913(.A(G208), .ZN(new_n1228_));
  OAI21_X1  g0914(.A(new_n1098_), .B1(new_n371_), .B2(new_n1228_), .ZN(new_n1229_));
  XNOR2_X1  g0915(.A(new_n1227_), .B(new_n1229_), .ZN(new_n1230_));
  NAND3_X1  g0916(.A1(new_n1224_), .A2(new_n1225_), .A3(new_n1230_), .ZN(new_n1231_));
  INV_X1    g0917(.A(new_n1225_), .ZN(new_n1232_));
  INV_X1    g0918(.A(new_n1230_), .ZN(new_n1233_));
  NAND3_X1  g0919(.A1(new_n1224_), .A2(new_n1232_), .A3(new_n1233_), .ZN(new_n1234_));
  NAND3_X1  g0920(.A1(new_n1223_), .A2(new_n1225_), .A3(new_n1233_), .ZN(new_n1235_));
  NAND3_X1  g0921(.A1(new_n1223_), .A2(new_n1232_), .A3(new_n1230_), .ZN(new_n1236_));
  NAND4_X1  g0922(.A1(new_n1231_), .A2(new_n1234_), .A3(new_n1235_), .A4(new_n1236_), .ZN(new_n1237_));
  XNOR2_X1  g0923(.A(new_n718_), .B(new_n712_), .ZN(new_n1238_));
  XOR2_X1   g0924(.A(new_n702_), .B(new_n707_), .Z(new_n1239_));
  XNOR2_X1  g0925(.A(new_n1238_), .B(new_n1239_), .ZN(new_n1240_));
  XNOR2_X1  g0926(.A(new_n1237_), .B(new_n1240_), .ZN(new_n1241_));
  XOR2_X1   g0927(.A(new_n871_), .B(new_n860_), .Z(new_n1242_));
  INV_X1    g0928(.A(new_n1242_), .ZN(new_n1243_));
  XNOR2_X1  g0929(.A(new_n854_), .B(new_n850_), .ZN(new_n1244_));
  INV_X1    g0930(.A(G197), .ZN(new_n1245_));
  OAI21_X1  g0931(.A(new_n1117_), .B1(new_n371_), .B2(new_n1245_), .ZN(new_n1246_));
  XNOR2_X1  g0932(.A(new_n867_), .B(new_n1246_), .ZN(new_n1247_));
  NAND3_X1  g0933(.A1(new_n1243_), .A2(new_n1244_), .A3(new_n1247_), .ZN(new_n1248_));
  INV_X1    g0934(.A(new_n1244_), .ZN(new_n1249_));
  INV_X1    g0935(.A(new_n1247_), .ZN(new_n1250_));
  NAND3_X1  g0936(.A1(new_n1243_), .A2(new_n1249_), .A3(new_n1250_), .ZN(new_n1251_));
  NAND3_X1  g0937(.A1(new_n1242_), .A2(new_n1244_), .A3(new_n1250_), .ZN(new_n1252_));
  NAND3_X1  g0938(.A1(new_n1242_), .A2(new_n1249_), .A3(new_n1247_), .ZN(new_n1253_));
  NAND4_X1  g0939(.A1(new_n1248_), .A2(new_n1251_), .A3(new_n1252_), .A4(new_n1253_), .ZN(new_n1254_));
  XNOR2_X1  g0940(.A(new_n877_), .B(new_n887_), .ZN(new_n1255_));
  XOR2_X1   g0941(.A(new_n882_), .B(new_n892_), .Z(new_n1256_));
  XNOR2_X1  g0942(.A(new_n1255_), .B(new_n1256_), .ZN(new_n1257_));
  XNOR2_X1  g0943(.A(new_n1254_), .B(new_n1257_), .ZN(new_n1258_));
  XNOR2_X1  g0944(.A(new_n772_), .B(new_n766_), .ZN(new_n1259_));
  INV_X1    g0945(.A(new_n1259_), .ZN(new_n1260_));
  XNOR2_X1  g0946(.A(new_n783_), .B(new_n778_), .ZN(new_n1261_));
  NOR3_X1   g0947(.A1(new_n377_), .A2(new_n371_), .A3(G170), .ZN(new_n1262_));
  NAND3_X1  g0948(.A1(new_n1260_), .A2(new_n1261_), .A3(new_n1262_), .ZN(new_n1263_));
  INV_X1    g0949(.A(new_n1261_), .ZN(new_n1264_));
  INV_X1    g0950(.A(new_n1262_), .ZN(new_n1265_));
  NAND3_X1  g0951(.A1(new_n1260_), .A2(new_n1264_), .A3(new_n1265_), .ZN(new_n1266_));
  NAND3_X1  g0952(.A1(new_n1259_), .A2(new_n1261_), .A3(new_n1265_), .ZN(new_n1267_));
  NAND3_X1  g0953(.A1(new_n1264_), .A2(new_n1259_), .A3(new_n1262_), .ZN(new_n1268_));
  NAND4_X1  g0954(.A1(new_n1263_), .A2(new_n1266_), .A3(new_n1267_), .A4(new_n1268_), .ZN(new_n1269_));
  OAI21_X1  g0955(.A(new_n383_), .B1(new_n371_), .B2(G165), .ZN(new_n1270_));
  OAI21_X1  g0956(.A(new_n383_), .B1(new_n371_), .B2(G164), .ZN(new_n1271_));
  XNOR2_X1  g0957(.A(new_n1270_), .B(new_n1271_), .ZN(new_n1272_));
  XNOR2_X1  g0958(.A(new_n1269_), .B(new_n1272_), .ZN(new_n1273_));
  NAND4_X1  g0959(.A1(new_n1222_), .A2(new_n1241_), .A3(new_n1258_), .A4(new_n1273_), .ZN(G416));
  INV_X1    g0960(.A(new_n929_), .ZN(new_n1275_));
  NAND3_X1  g0961(.A1(new_n764_), .A2(new_n845_), .A3(new_n899_), .ZN(new_n1276_));
  NOR2_X1   g0962(.A1(new_n917_), .A2(new_n927_), .ZN(new_n1277_));
  NAND2_X1  g0963(.A1(new_n963_), .A2(new_n845_), .ZN(new_n1278_));
  NAND4_X1  g0964(.A1(new_n899_), .A2(new_n904_), .A3(G89), .A4(new_n845_), .ZN(new_n1279_));
  NAND4_X1  g0965(.A1(new_n1276_), .A2(new_n1277_), .A3(new_n1278_), .A4(new_n1279_), .ZN(new_n1280_));
  AOI21_X1  g0966(.A(new_n942_), .B1(new_n1280_), .B2(new_n788_), .ZN(new_n1281_));
  INV_X1    g0967(.A(new_n795_), .ZN(new_n1282_));
  OAI21_X1  g0968(.A(new_n1275_), .B1(new_n1281_), .B2(new_n1282_), .ZN(G249));
  AOI21_X1  g0969(.A(new_n607_), .B1(new_n533_), .B2(new_n548_), .ZN(new_n1284_));
  NAND3_X1  g0970(.A1(new_n613_), .A2(new_n608_), .A3(G4526), .ZN(new_n1285_));
  NAND3_X1  g0971(.A1(new_n687_), .A2(new_n697_), .A3(new_n1285_), .ZN(new_n1286_));
  NOR2_X1   g0972(.A1(new_n1284_), .A2(new_n1286_), .ZN(new_n1287_));
  XNOR2_X1  g0973(.A(new_n1287_), .B(new_n459_), .ZN(G295));
  NAND2_X1  g0974(.A1(new_n533_), .A2(new_n548_), .ZN(new_n1289_));
  NAND3_X1  g0975(.A1(new_n1289_), .A2(new_n462_), .A3(new_n608_), .ZN(new_n1290_));
  NAND2_X1  g0976(.A1(new_n698_), .A2(new_n462_), .ZN(new_n1291_));
  NAND4_X1  g0977(.A1(new_n613_), .A2(new_n608_), .A3(G4526), .A4(new_n462_), .ZN(new_n1292_));
  NAND4_X1  g0978(.A1(new_n1290_), .A2(new_n643_), .A3(new_n1291_), .A4(new_n1292_), .ZN(new_n1293_));
  XNOR2_X1  g0979(.A(new_n1293_), .B(new_n398_), .ZN(G324));
  INV_X1    g0980(.A(G89), .ZN(new_n1295_));
  NOR2_X1   g0981(.A1(new_n903_), .A2(new_n1295_), .ZN(new_n1296_));
  NOR3_X1   g0982(.A1(new_n759_), .A2(new_n760_), .A3(new_n1296_), .ZN(new_n1297_));
  OAI21_X1  g0983(.A(new_n725_), .B1(new_n1297_), .B2(new_n763_), .ZN(new_n1298_));
  AOI21_X1  g0984(.A(new_n955_), .B1(new_n1298_), .B2(new_n875_), .ZN(new_n1299_));
  OAI21_X1  g0985(.A(new_n962_), .B1(new_n1299_), .B2(new_n896_), .ZN(G252));
  NOR2_X1   g0986(.A1(new_n1001_), .A2(new_n627_), .ZN(new_n1301_));
  NAND2_X1  g0987(.A1(new_n1005_), .A2(new_n991_), .ZN(new_n1302_));
  NAND4_X1  g0988(.A1(new_n998_), .A2(G4526), .A3(new_n991_), .A4(new_n979_), .ZN(new_n1303_));
  NAND3_X1  g0989(.A1(new_n969_), .A2(new_n991_), .A3(new_n979_), .ZN(new_n1304_));
  NAND4_X1  g0990(.A1(new_n1301_), .A2(new_n1302_), .A3(new_n1303_), .A4(new_n1304_), .ZN(new_n1305_));
  AOI21_X1  g0991(.A(new_n667_), .B1(new_n1305_), .B2(new_n983_), .ZN(new_n1306_));
  OAI21_X1  g0992(.A(new_n645_), .B1(new_n1306_), .B2(new_n985_), .ZN(G276));
  INV_X1    g0993(.A(new_n1287_), .ZN(new_n1308_));
  INV_X1    g0994(.A(new_n438_), .ZN(new_n1309_));
  AOI21_X1  g0995(.A(new_n437_), .B1(new_n804_), .B2(new_n433_), .ZN(new_n1310_));
  NOR2_X1   g0996(.A1(new_n1309_), .A2(new_n1310_), .ZN(new_n1311_));
  NOR3_X1   g0997(.A1(new_n455_), .A2(new_n1311_), .A3(new_n989_), .ZN(new_n1312_));
  NAND3_X1  g0998(.A1(new_n1308_), .A2(new_n459_), .A3(new_n1312_), .ZN(new_n1313_));
  NAND4_X1  g0999(.A1(new_n454_), .A2(new_n439_), .A3(new_n446_), .A4(new_n628_), .ZN(new_n1314_));
  AND2_X1   g1000(.A1(new_n1313_), .A2(new_n1314_), .ZN(new_n1315_));
  NAND3_X1  g1001(.A1(new_n454_), .A2(new_n439_), .A3(new_n637_), .ZN(new_n1316_));
  NAND4_X1  g1002(.A1(new_n1315_), .A2(new_n640_), .A3(new_n633_), .A4(new_n1316_), .ZN(new_n1317_));
  XNOR2_X1  g1003(.A(new_n1317_), .B(new_n431_), .ZN(G310));
  NAND4_X1  g1004(.A1(new_n1308_), .A2(new_n439_), .A3(new_n446_), .A4(new_n459_), .ZN(new_n1319_));
  NAND2_X1  g1005(.A1(new_n435_), .A2(new_n437_), .ZN(new_n1320_));
  OAI21_X1  g1006(.A(new_n637_), .B1(new_n1309_), .B2(new_n1310_), .ZN(new_n1321_));
  NAND3_X1  g1007(.A1(new_n439_), .A2(new_n446_), .A3(new_n628_), .ZN(new_n1322_));
  NAND4_X1  g1008(.A1(new_n1319_), .A2(new_n1320_), .A3(new_n1321_), .A4(new_n1322_), .ZN(new_n1323_));
  XNOR2_X1  g1009(.A(new_n1323_), .B(new_n455_), .ZN(G313));
  NAND3_X1  g1010(.A1(new_n1308_), .A2(new_n446_), .A3(new_n459_), .ZN(new_n1325_));
  INV_X1    g1011(.A(new_n637_), .ZN(new_n1326_));
  INV_X1    g1012(.A(new_n445_), .ZN(new_n1327_));
  AOI21_X1  g1013(.A(new_n444_), .B1(new_n636_), .B2(new_n440_), .ZN(new_n1328_));
  OAI21_X1  g1014(.A(new_n628_), .B1(new_n1327_), .B2(new_n1328_), .ZN(new_n1329_));
  NAND3_X1  g1015(.A1(new_n1325_), .A2(new_n1326_), .A3(new_n1329_), .ZN(new_n1330_));
  XNOR2_X1  g1016(.A(new_n1330_), .B(new_n1311_), .ZN(G316));
  OAI21_X1  g1017(.A(new_n629_), .B1(new_n1287_), .B2(new_n460_), .ZN(new_n1332_));
  XNOR2_X1  g1018(.A(new_n1332_), .B(new_n989_), .ZN(G319));
  INV_X1    g1019(.A(new_n387_), .ZN(new_n1334_));
  AOI21_X1  g1020(.A(G106), .B1(new_n652_), .B2(new_n383_), .ZN(new_n1335_));
  NOR2_X1   g1021(.A1(new_n1334_), .A2(new_n1335_), .ZN(new_n1336_));
  NOR3_X1   g1022(.A1(new_n405_), .A2(new_n982_), .A3(new_n1336_), .ZN(new_n1337_));
  NAND3_X1  g1023(.A1(new_n1293_), .A2(new_n397_), .A3(new_n1337_), .ZN(new_n1338_));
  NAND3_X1  g1024(.A1(new_n404_), .A2(new_n388_), .A3(new_n661_), .ZN(new_n1339_));
  INV_X1    g1025(.A(new_n647_), .ZN(new_n1340_));
  NAND4_X1  g1026(.A1(new_n404_), .A2(new_n388_), .A3(new_n393_), .A4(new_n1340_), .ZN(new_n1341_));
  NAND4_X1  g1027(.A1(new_n1338_), .A2(new_n664_), .A3(new_n1339_), .A4(new_n1341_), .ZN(new_n1342_));
  NOR2_X1   g1028(.A1(new_n1342_), .A2(new_n656_), .ZN(new_n1343_));
  XNOR2_X1  g1029(.A(new_n1343_), .B(new_n382_), .ZN(G327));
  NAND4_X1  g1030(.A1(new_n1293_), .A2(new_n397_), .A3(new_n388_), .A4(new_n393_), .ZN(new_n1345_));
  OAI21_X1  g1031(.A(new_n661_), .B1(new_n1334_), .B2(new_n1335_), .ZN(new_n1346_));
  AOI21_X1  g1032(.A(new_n647_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n1347_));
  NAND2_X1  g1033(.A1(new_n1347_), .A2(new_n388_), .ZN(new_n1348_));
  NAND4_X1  g1034(.A1(new_n1345_), .A2(new_n653_), .A3(new_n1346_), .A4(new_n1348_), .ZN(new_n1349_));
  XNOR2_X1  g1035(.A(new_n1349_), .B(new_n405_), .ZN(G330));
  NAND3_X1  g1036(.A1(new_n1293_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n1351_));
  INV_X1    g1037(.A(new_n392_), .ZN(new_n1352_));
  AOI21_X1  g1038(.A(G1469), .B1(new_n659_), .B2(new_n383_), .ZN(new_n1353_));
  OAI21_X1  g1039(.A(new_n1340_), .B1(new_n1352_), .B2(new_n1353_), .ZN(new_n1354_));
  NAND3_X1  g1040(.A1(new_n1351_), .A2(new_n660_), .A3(new_n1354_), .ZN(new_n1355_));
  XNOR2_X1  g1041(.A(new_n1355_), .B(new_n1336_), .ZN(G333));
  AOI21_X1  g1042(.A(new_n1340_), .B1(new_n1293_), .B2(new_n397_), .ZN(new_n1357_));
  XNOR2_X1  g1043(.A(new_n1357_), .B(new_n393_), .ZN(G336));
  NOR3_X1   g1044(.A1(G416), .A2(G412), .A3(G414), .ZN(new_n1359_));
  NOR2_X1   g1045(.A1(G408), .A2(G410), .ZN(new_n1360_));
  NOR2_X1   g1046(.A1(G404), .A2(G406), .ZN(new_n1361_));
  NAND3_X1  g1047(.A1(new_n1359_), .A2(new_n1360_), .A3(new_n1361_), .ZN(G418));
  NAND2_X1  g1048(.A1(new_n1293_), .A2(new_n406_), .ZN(new_n1363_));
  NAND2_X1  g1049(.A1(new_n1363_), .A2(new_n666_), .ZN(new_n1364_));
  INV_X1    g1050(.A(new_n1364_), .ZN(new_n1365_));
  OAI21_X1  g1051(.A(new_n645_), .B1(new_n1365_), .B2(new_n985_), .ZN(G273));
  AOI21_X1  g1052(.A(new_n642_), .B1(new_n1308_), .B2(new_n461_), .ZN(new_n1367_));
  NAND3_X1  g1053(.A1(new_n619_), .A2(new_n620_), .A3(new_n626_), .ZN(new_n1368_));
  XNOR2_X1  g1054(.A(new_n1368_), .B(new_n426_), .ZN(new_n1369_));
  NAND2_X1  g1055(.A1(new_n1367_), .A2(new_n1369_), .ZN(new_n1370_));
  OAI211_X1 g1056(.A(new_n416_), .B(new_n423_), .C1(new_n616_), .C2(new_n615_), .ZN(new_n1371_));
  NAND3_X1  g1057(.A1(new_n1371_), .A2(new_n626_), .A3(new_n620_), .ZN(new_n1372_));
  INV_X1    g1058(.A(new_n426_), .ZN(new_n1373_));
  XNOR2_X1  g1059(.A(new_n1372_), .B(new_n1373_), .ZN(new_n1374_));
  OAI21_X1  g1060(.A(new_n1370_), .B1(new_n1367_), .B2(new_n1374_), .ZN(G298));
  NAND2_X1  g1061(.A1(new_n423_), .A2(new_n618_), .ZN(new_n1376_));
  NAND2_X1  g1062(.A1(new_n419_), .A2(new_n421_), .ZN(new_n1377_));
  NAND2_X1  g1063(.A1(new_n1376_), .A2(new_n1377_), .ZN(new_n1378_));
  XNOR2_X1  g1064(.A(new_n1378_), .B(new_n417_), .ZN(new_n1379_));
  NAND2_X1  g1065(.A1(new_n1367_), .A2(new_n1379_), .ZN(new_n1380_));
  OAI211_X1 g1066(.A(new_n1376_), .B(new_n1377_), .C1(new_n424_), .C2(new_n428_), .ZN(new_n1381_));
  XNOR2_X1  g1067(.A(new_n1381_), .B(new_n416_), .ZN(new_n1382_));
  OAI21_X1  g1068(.A(new_n1380_), .B1(new_n1367_), .B2(new_n1382_), .ZN(G301));
  XNOR2_X1  g1069(.A(new_n423_), .B(new_n617_), .ZN(new_n1384_));
  NAND2_X1  g1070(.A1(new_n1367_), .A2(new_n1384_), .ZN(new_n1385_));
  NAND2_X1  g1071(.A1(new_n427_), .A2(G2239), .ZN(new_n1386_));
  XNOR2_X1  g1072(.A(new_n423_), .B(new_n1386_), .ZN(new_n1387_));
  OAI21_X1  g1073(.A(new_n1385_), .B1(new_n1367_), .B2(new_n1387_), .ZN(G304));
  INV_X1    g1074(.A(new_n428_), .ZN(new_n1389_));
  XNOR2_X1  g1075(.A(new_n1367_), .B(new_n1389_), .ZN(G307));
  INV_X1    g1076(.A(new_n532_), .ZN(new_n1391_));
  OAI21_X1  g1077(.A(new_n548_), .B1(new_n1035_), .B2(new_n1391_), .ZN(new_n1392_));
  XNOR2_X1  g1078(.A(new_n1392_), .B(new_n605_), .ZN(G344));
  NOR2_X1   g1079(.A1(new_n407_), .A2(G38), .ZN(new_n1394_));
  XOR2_X1   g1080(.A(new_n410_), .B(new_n1394_), .Z(new_n1395_));
  NAND2_X1  g1081(.A1(new_n1364_), .A2(new_n1395_), .ZN(new_n1396_));
  NAND2_X1  g1082(.A1(new_n407_), .A2(G38), .ZN(new_n1397_));
  XNOR2_X1  g1083(.A(new_n410_), .B(new_n1397_), .ZN(new_n1398_));
  OAI21_X1  g1084(.A(new_n1396_), .B1(new_n1364_), .B2(new_n1398_), .ZN(G422));
  OAI21_X1  g1085(.A(new_n1396_), .B1(new_n1364_), .B2(new_n1398_), .ZN(G469));
  XNOR2_X1  g1086(.A(new_n1364_), .B(new_n408_), .ZN(G419));
  XNOR2_X1  g1087(.A(new_n1364_), .B(new_n408_), .ZN(G471));
  INV_X1    g1088(.A(new_n599_), .ZN(new_n1403_));
  NOR3_X1   g1089(.A1(new_n669_), .A2(new_n973_), .A3(new_n1403_), .ZN(new_n1404_));
  NAND3_X1  g1090(.A1(new_n1392_), .A2(new_n604_), .A3(new_n1404_), .ZN(new_n1405_));
  NAND3_X1  g1091(.A1(new_n585_), .A2(new_n592_), .A3(new_n680_), .ZN(new_n1406_));
  NAND4_X1  g1092(.A1(new_n585_), .A2(new_n592_), .A3(new_n599_), .A4(new_n670_), .ZN(new_n1407_));
  NAND4_X1  g1093(.A1(new_n1405_), .A2(new_n684_), .A3(new_n1406_), .A4(new_n1407_), .ZN(new_n1408_));
  NOR2_X1   g1094(.A1(new_n1408_), .A2(new_n677_), .ZN(new_n1409_));
  XNOR2_X1  g1095(.A(new_n1409_), .B(new_n578_), .ZN(G359));
  NAND4_X1  g1096(.A1(new_n1392_), .A2(new_n592_), .A3(new_n599_), .A4(new_n604_), .ZN(new_n1411_));
  NAND2_X1  g1097(.A1(new_n588_), .A2(new_n590_), .ZN(new_n1412_));
  OAI21_X1  g1098(.A(new_n680_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n1413_));
  NAND3_X1  g1099(.A1(new_n592_), .A2(new_n599_), .A3(new_n670_), .ZN(new_n1414_));
  NAND4_X1  g1100(.A1(new_n1411_), .A2(new_n1412_), .A3(new_n1413_), .A4(new_n1414_), .ZN(new_n1415_));
  XNOR2_X1  g1101(.A(new_n1415_), .B(new_n669_), .ZN(G362));
  NAND3_X1  g1102(.A1(new_n1392_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n1417_));
  INV_X1    g1103(.A(new_n680_), .ZN(new_n1418_));
  INV_X1    g1104(.A(new_n598_), .ZN(new_n1419_));
  AOI21_X1  g1105(.A(new_n597_), .B1(new_n679_), .B2(new_n593_), .ZN(new_n1420_));
  OAI21_X1  g1106(.A(new_n670_), .B1(new_n1419_), .B2(new_n1420_), .ZN(new_n1421_));
  NAND3_X1  g1107(.A1(new_n1417_), .A2(new_n1418_), .A3(new_n1421_), .ZN(new_n1422_));
  XNOR2_X1  g1108(.A(new_n1422_), .B(new_n973_), .ZN(G365));
  AOI21_X1  g1109(.A(new_n670_), .B1(new_n1392_), .B2(new_n604_), .ZN(new_n1424_));
  XNOR2_X1  g1110(.A(new_n1424_), .B(new_n599_), .ZN(G368));
  AOI21_X1  g1111(.A(new_n686_), .B1(new_n1392_), .B2(new_n606_), .ZN(new_n1426_));
  NAND3_X1  g1112(.A1(new_n693_), .A2(new_n689_), .A3(new_n695_), .ZN(new_n1427_));
  XNOR2_X1  g1113(.A(new_n1427_), .B(new_n568_), .ZN(new_n1428_));
  NAND2_X1  g1114(.A1(new_n1426_), .A2(new_n1428_), .ZN(new_n1429_));
  OAI211_X1 g1115(.A(new_n553_), .B(new_n562_), .C1(new_n572_), .C2(new_n571_), .ZN(new_n1430_));
  NAND3_X1  g1116(.A1(new_n1430_), .A2(new_n689_), .A3(new_n695_), .ZN(new_n1431_));
  XNOR2_X1  g1117(.A(new_n1431_), .B(new_n976_), .ZN(new_n1432_));
  OAI21_X1  g1118(.A(new_n1429_), .B1(new_n1426_), .B2(new_n1432_), .ZN(G347));
  NAND2_X1  g1119(.A1(new_n562_), .A2(new_n692_), .ZN(new_n1434_));
  INV_X1    g1120(.A(new_n694_), .ZN(new_n1435_));
  NAND2_X1  g1121(.A1(new_n1434_), .A2(new_n1435_), .ZN(new_n1436_));
  XNOR2_X1  g1122(.A(new_n1436_), .B(new_n554_), .ZN(new_n1437_));
  NAND2_X1  g1123(.A1(new_n1426_), .A2(new_n1437_), .ZN(new_n1438_));
  OAI211_X1 g1124(.A(new_n1434_), .B(new_n1435_), .C1(new_n563_), .C2(new_n573_), .ZN(new_n1439_));
  XNOR2_X1  g1125(.A(new_n1439_), .B(new_n553_), .ZN(new_n1440_));
  OAI21_X1  g1126(.A(new_n1438_), .B1(new_n1426_), .B2(new_n1440_), .ZN(G350));
  INV_X1    g1127(.A(new_n692_), .ZN(new_n1442_));
  XNOR2_X1  g1128(.A(new_n1442_), .B(new_n562_), .ZN(new_n1443_));
  NAND2_X1  g1129(.A1(new_n1426_), .A2(new_n1443_), .ZN(new_n1444_));
  NAND2_X1  g1130(.A1(new_n691_), .A2(G4420), .ZN(new_n1445_));
  XNOR2_X1  g1131(.A(new_n562_), .B(new_n1445_), .ZN(new_n1446_));
  OAI21_X1  g1132(.A(new_n1444_), .B1(new_n1426_), .B2(new_n1446_), .ZN(G353));
  XNOR2_X1  g1133(.A(new_n1426_), .B(new_n977_), .ZN(G356));
  AND2_X1   g1134(.A1(new_n1004_), .A2(new_n697_), .ZN(new_n1449_));
  NAND3_X1  g1135(.A1(new_n998_), .A2(G4526), .A3(new_n979_), .ZN(new_n1450_));
  OAI211_X1 g1136(.A(new_n1449_), .B(new_n1450_), .C1(new_n970_), .C2(new_n980_), .ZN(new_n1451_));
  INV_X1    g1137(.A(new_n1451_), .ZN(new_n1452_));
  NAND4_X1  g1138(.A1(new_n459_), .A2(new_n454_), .A3(new_n439_), .A4(new_n446_), .ZN(new_n1453_));
  NAND4_X1  g1139(.A1(new_n1453_), .A2(new_n1314_), .A3(new_n640_), .A4(new_n1316_), .ZN(new_n1454_));
  NOR2_X1   g1140(.A1(new_n1454_), .A2(new_n634_), .ZN(new_n1455_));
  INV_X1    g1141(.A(G2211), .ZN(new_n1456_));
  OAI211_X1 g1142(.A(new_n439_), .B(new_n446_), .C1(new_n1456_), .C2(new_n458_), .ZN(new_n1457_));
  NAND3_X1  g1143(.A1(new_n1457_), .A2(new_n1320_), .A3(new_n1321_), .ZN(new_n1458_));
  INV_X1    g1144(.A(new_n458_), .ZN(new_n1459_));
  NAND2_X1  g1145(.A1(new_n1459_), .A2(G2211), .ZN(new_n1460_));
  NAND2_X1  g1146(.A1(new_n1458_), .A2(new_n1460_), .ZN(new_n1461_));
  NAND2_X1  g1147(.A1(new_n1329_), .A2(new_n1326_), .ZN(new_n1462_));
  INV_X1    g1148(.A(new_n1462_), .ZN(new_n1463_));
  OAI21_X1  g1149(.A(new_n1463_), .B1(new_n989_), .B2(new_n460_), .ZN(new_n1464_));
  INV_X1    g1150(.A(new_n1460_), .ZN(new_n1465_));
  NAND4_X1  g1151(.A1(new_n1457_), .A2(new_n1320_), .A3(new_n1321_), .A4(new_n1465_), .ZN(new_n1466_));
  AND3_X1   g1152(.A1(new_n1461_), .A2(new_n1464_), .A3(new_n1466_), .ZN(new_n1467_));
  AOI21_X1  g1153(.A(new_n1464_), .B1(new_n1461_), .B2(new_n1466_), .ZN(new_n1468_));
  OAI21_X1  g1154(.A(new_n1455_), .B1(new_n1467_), .B2(new_n1468_), .ZN(new_n1469_));
  NAND2_X1  g1155(.A1(new_n1461_), .A2(new_n1466_), .ZN(new_n1470_));
  INV_X1    g1156(.A(new_n1464_), .ZN(new_n1471_));
  NAND2_X1  g1157(.A1(new_n1470_), .A2(new_n1471_), .ZN(new_n1472_));
  OR2_X1    g1158(.A1(new_n1454_), .A2(new_n634_), .ZN(new_n1473_));
  NAND3_X1  g1159(.A1(new_n1461_), .A2(new_n1464_), .A3(new_n1466_), .ZN(new_n1474_));
  NAND3_X1  g1160(.A1(new_n1472_), .A2(new_n1473_), .A3(new_n1474_), .ZN(new_n1475_));
  AND3_X1   g1161(.A1(new_n1469_), .A2(new_n1475_), .A3(new_n459_), .ZN(new_n1476_));
  AOI21_X1  g1162(.A(new_n459_), .B1(new_n1469_), .B2(new_n1475_), .ZN(new_n1477_));
  OAI21_X1  g1163(.A(new_n989_), .B1(new_n1476_), .B2(new_n1477_), .ZN(new_n1478_));
  NOR3_X1   g1164(.A1(new_n1467_), .A2(new_n1468_), .A3(new_n1455_), .ZN(new_n1479_));
  AOI21_X1  g1165(.A(new_n1473_), .B1(new_n1472_), .B2(new_n1474_), .ZN(new_n1480_));
  OAI21_X1  g1166(.A(new_n460_), .B1(new_n1479_), .B2(new_n1480_), .ZN(new_n1481_));
  NAND3_X1  g1167(.A1(new_n1469_), .A2(new_n1475_), .A3(new_n459_), .ZN(new_n1482_));
  NAND3_X1  g1168(.A1(new_n1481_), .A2(new_n446_), .A3(new_n1482_), .ZN(new_n1483_));
  AND3_X1   g1169(.A1(new_n1478_), .A2(new_n432_), .A3(new_n1483_), .ZN(new_n1484_));
  AOI21_X1  g1170(.A(new_n432_), .B1(new_n1478_), .B2(new_n1483_), .ZN(new_n1485_));
  NOR3_X1   g1171(.A1(new_n1484_), .A2(new_n1485_), .A3(new_n1311_), .ZN(new_n1486_));
  NOR3_X1   g1172(.A1(new_n1476_), .A2(new_n1477_), .A3(new_n989_), .ZN(new_n1487_));
  AOI21_X1  g1173(.A(new_n446_), .B1(new_n1481_), .B2(new_n1482_), .ZN(new_n1488_));
  OAI21_X1  g1174(.A(new_n431_), .B1(new_n1487_), .B2(new_n1488_), .ZN(new_n1489_));
  NAND3_X1  g1175(.A1(new_n1478_), .A2(new_n1483_), .A3(new_n432_), .ZN(new_n1490_));
  AOI21_X1  g1176(.A(new_n439_), .B1(new_n1489_), .B2(new_n1490_), .ZN(new_n1491_));
  OAI21_X1  g1177(.A(new_n455_), .B1(new_n1486_), .B2(new_n1491_), .ZN(new_n1492_));
  OAI21_X1  g1178(.A(new_n1311_), .B1(new_n1484_), .B2(new_n1485_), .ZN(new_n1493_));
  NAND3_X1  g1179(.A1(new_n1489_), .A2(new_n439_), .A3(new_n1490_), .ZN(new_n1494_));
  NAND3_X1  g1180(.A1(new_n1493_), .A2(new_n454_), .A3(new_n1494_), .ZN(new_n1495_));
  AOI21_X1  g1181(.A(new_n1452_), .B1(new_n1492_), .B2(new_n1495_), .ZN(new_n1496_));
  NAND4_X1  g1182(.A1(new_n1314_), .A2(new_n633_), .A3(new_n1316_), .A4(new_n640_), .ZN(new_n1497_));
  OAI211_X1 g1183(.A(new_n1320_), .B(new_n1321_), .C1(new_n1329_), .C2(new_n1311_), .ZN(new_n1498_));
  NAND2_X1  g1184(.A1(new_n1498_), .A2(new_n628_), .ZN(new_n1499_));
  NAND4_X1  g1185(.A1(new_n1322_), .A2(new_n1320_), .A3(new_n629_), .A4(new_n1321_), .ZN(new_n1500_));
  AND3_X1   g1186(.A1(new_n1499_), .A2(new_n1463_), .A3(new_n1500_), .ZN(new_n1501_));
  AOI21_X1  g1187(.A(new_n1463_), .B1(new_n1499_), .B2(new_n1500_), .ZN(new_n1502_));
  OAI21_X1  g1188(.A(new_n1497_), .B1(new_n1501_), .B2(new_n1502_), .ZN(new_n1503_));
  NAND2_X1  g1189(.A1(new_n1499_), .A2(new_n1500_), .ZN(new_n1504_));
  NAND2_X1  g1190(.A1(new_n1504_), .A2(new_n1462_), .ZN(new_n1505_));
  INV_X1    g1191(.A(new_n1497_), .ZN(new_n1506_));
  NAND3_X1  g1192(.A1(new_n1499_), .A2(new_n1463_), .A3(new_n1500_), .ZN(new_n1507_));
  NAND3_X1  g1193(.A1(new_n1505_), .A2(new_n1506_), .A3(new_n1507_), .ZN(new_n1508_));
  AND3_X1   g1194(.A1(new_n1503_), .A2(new_n1508_), .A3(new_n459_), .ZN(new_n1509_));
  AOI21_X1  g1195(.A(new_n459_), .B1(new_n1503_), .B2(new_n1508_), .ZN(new_n1510_));
  OAI21_X1  g1196(.A(new_n989_), .B1(new_n1509_), .B2(new_n1510_), .ZN(new_n1511_));
  NOR3_X1   g1197(.A1(new_n1501_), .A2(new_n1502_), .A3(new_n1497_), .ZN(new_n1512_));
  AOI21_X1  g1198(.A(new_n1506_), .B1(new_n1505_), .B2(new_n1507_), .ZN(new_n1513_));
  OAI21_X1  g1199(.A(new_n460_), .B1(new_n1512_), .B2(new_n1513_), .ZN(new_n1514_));
  NAND3_X1  g1200(.A1(new_n1503_), .A2(new_n1508_), .A3(new_n459_), .ZN(new_n1515_));
  NAND3_X1  g1201(.A1(new_n1514_), .A2(new_n446_), .A3(new_n1515_), .ZN(new_n1516_));
  AND3_X1   g1202(.A1(new_n1511_), .A2(new_n432_), .A3(new_n1516_), .ZN(new_n1517_));
  AOI21_X1  g1203(.A(new_n432_), .B1(new_n1511_), .B2(new_n1516_), .ZN(new_n1518_));
  OAI21_X1  g1204(.A(new_n1311_), .B1(new_n1517_), .B2(new_n1518_), .ZN(new_n1519_));
  NOR3_X1   g1205(.A1(new_n1509_), .A2(new_n1510_), .A3(new_n989_), .ZN(new_n1520_));
  AOI21_X1  g1206(.A(new_n446_), .B1(new_n1514_), .B2(new_n1515_), .ZN(new_n1521_));
  OAI21_X1  g1207(.A(new_n431_), .B1(new_n1520_), .B2(new_n1521_), .ZN(new_n1522_));
  NAND3_X1  g1208(.A1(new_n1511_), .A2(new_n1516_), .A3(new_n432_), .ZN(new_n1523_));
  NAND3_X1  g1209(.A1(new_n1522_), .A2(new_n439_), .A3(new_n1523_), .ZN(new_n1524_));
  AND3_X1   g1210(.A1(new_n1519_), .A2(new_n454_), .A3(new_n1524_), .ZN(new_n1525_));
  AOI21_X1  g1211(.A(new_n454_), .B1(new_n1519_), .B2(new_n1524_), .ZN(new_n1526_));
  NOR3_X1   g1212(.A1(new_n1525_), .A2(new_n1526_), .A3(new_n1451_), .ZN(new_n1527_));
  OAI22_X1  g1213(.A1(new_n616_), .A2(new_n615_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n1528_));
  OAI211_X1 g1214(.A(G2239), .B(new_n427_), .C1(new_n418_), .C2(G2247), .ZN(new_n1529_));
  NAND2_X1  g1215(.A1(new_n1528_), .A2(new_n1529_), .ZN(new_n1530_));
  INV_X1    g1216(.A(new_n1530_), .ZN(new_n1531_));
  NAND2_X1  g1217(.A1(new_n1372_), .A2(new_n1531_), .ZN(new_n1532_));
  NAND4_X1  g1218(.A1(new_n1371_), .A2(new_n626_), .A3(new_n620_), .A4(new_n1530_), .ZN(new_n1533_));
  AOI21_X1  g1219(.A(new_n1389_), .B1(new_n1532_), .B2(new_n1533_), .ZN(new_n1534_));
  INV_X1    g1220(.A(new_n1534_), .ZN(new_n1535_));
  NAND3_X1  g1221(.A1(new_n1532_), .A2(new_n1389_), .A3(new_n1533_), .ZN(new_n1536_));
  AOI21_X1  g1222(.A(new_n423_), .B1(new_n1535_), .B2(new_n1536_), .ZN(new_n1537_));
  INV_X1    g1223(.A(new_n1536_), .ZN(new_n1538_));
  NOR3_X1   g1224(.A1(new_n1538_), .A2(new_n424_), .A3(new_n1534_), .ZN(new_n1539_));
  OAI21_X1  g1225(.A(new_n426_), .B1(new_n1537_), .B2(new_n1539_), .ZN(new_n1540_));
  OAI21_X1  g1226(.A(new_n424_), .B1(new_n1538_), .B2(new_n1534_), .ZN(new_n1541_));
  NAND3_X1  g1227(.A1(new_n1535_), .A2(new_n423_), .A3(new_n1536_), .ZN(new_n1542_));
  NAND3_X1  g1228(.A1(new_n1541_), .A2(new_n1542_), .A3(new_n1373_), .ZN(new_n1543_));
  AND3_X1   g1229(.A1(new_n1540_), .A2(new_n416_), .A3(new_n1543_), .ZN(new_n1544_));
  AOI21_X1  g1230(.A(new_n416_), .B1(new_n1540_), .B2(new_n1543_), .ZN(new_n1545_));
  OAI211_X1 g1231(.A(new_n642_), .B(new_n1452_), .C1(new_n1544_), .C2(new_n1545_), .ZN(new_n1546_));
  NOR2_X1   g1232(.A1(new_n642_), .A2(new_n990_), .ZN(new_n1547_));
  INV_X1    g1233(.A(new_n1547_), .ZN(new_n1548_));
  OAI211_X1 g1234(.A(new_n1451_), .B(new_n1548_), .C1(new_n1544_), .C2(new_n1545_), .ZN(new_n1549_));
  INV_X1    g1235(.A(new_n642_), .ZN(new_n1550_));
  NAND3_X1  g1236(.A1(new_n416_), .A2(new_n423_), .A3(new_n618_), .ZN(new_n1551_));
  NAND3_X1  g1237(.A1(new_n620_), .A2(new_n1551_), .A3(new_n626_), .ZN(new_n1552_));
  OAI21_X1  g1238(.A(new_n618_), .B1(new_n421_), .B2(new_n419_), .ZN(new_n1553_));
  OAI21_X1  g1239(.A(new_n617_), .B1(G2247), .B2(new_n418_), .ZN(new_n1554_));
  NAND2_X1  g1240(.A1(new_n1553_), .A2(new_n1554_), .ZN(new_n1555_));
  NAND2_X1  g1241(.A1(new_n1552_), .A2(new_n1555_), .ZN(new_n1556_));
  INV_X1    g1242(.A(new_n1555_), .ZN(new_n1557_));
  NAND4_X1  g1243(.A1(new_n1557_), .A2(new_n626_), .A3(new_n620_), .A4(new_n1551_), .ZN(new_n1558_));
  AOI21_X1  g1244(.A(new_n1389_), .B1(new_n1556_), .B2(new_n1558_), .ZN(new_n1559_));
  INV_X1    g1245(.A(new_n1559_), .ZN(new_n1560_));
  NAND3_X1  g1246(.A1(new_n1556_), .A2(new_n1558_), .A3(new_n1389_), .ZN(new_n1561_));
  AOI21_X1  g1247(.A(new_n423_), .B1(new_n1560_), .B2(new_n1561_), .ZN(new_n1562_));
  INV_X1    g1248(.A(new_n1561_), .ZN(new_n1563_));
  NOR3_X1   g1249(.A1(new_n1563_), .A2(new_n1559_), .A3(new_n424_), .ZN(new_n1564_));
  OAI21_X1  g1250(.A(new_n426_), .B1(new_n1562_), .B2(new_n1564_), .ZN(new_n1565_));
  NAND3_X1  g1251(.A1(new_n1560_), .A2(new_n423_), .A3(new_n1561_), .ZN(new_n1566_));
  OAI21_X1  g1252(.A(new_n424_), .B1(new_n1563_), .B2(new_n1559_), .ZN(new_n1567_));
  NAND3_X1  g1253(.A1(new_n1566_), .A2(new_n1567_), .A3(new_n1373_), .ZN(new_n1568_));
  AND3_X1   g1254(.A1(new_n1565_), .A2(new_n416_), .A3(new_n1568_), .ZN(new_n1569_));
  AOI21_X1  g1255(.A(new_n416_), .B1(new_n1565_), .B2(new_n1568_), .ZN(new_n1570_));
  OAI211_X1 g1256(.A(new_n1452_), .B(new_n1550_), .C1(new_n1569_), .C2(new_n1570_), .ZN(new_n1571_));
  OAI211_X1 g1257(.A(new_n1451_), .B(new_n1547_), .C1(new_n1569_), .C2(new_n1570_), .ZN(new_n1572_));
  AND4_X1   g1258(.A1(new_n1546_), .A2(new_n1549_), .A3(new_n1571_), .A4(new_n1572_), .ZN(new_n1573_));
  NOR3_X1   g1259(.A1(new_n1496_), .A2(new_n1527_), .A3(new_n1573_), .ZN(new_n1574_));
  NAND4_X1  g1260(.A1(new_n1546_), .A2(new_n1549_), .A3(new_n1571_), .A4(new_n1572_), .ZN(new_n1575_));
  AND3_X1   g1261(.A1(new_n1493_), .A2(new_n454_), .A3(new_n1494_), .ZN(new_n1576_));
  AOI21_X1  g1262(.A(new_n454_), .B1(new_n1493_), .B2(new_n1494_), .ZN(new_n1577_));
  OAI21_X1  g1263(.A(new_n1451_), .B1(new_n1576_), .B2(new_n1577_), .ZN(new_n1578_));
  INV_X1    g1264(.A(new_n1526_), .ZN(new_n1579_));
  NAND3_X1  g1265(.A1(new_n1519_), .A2(new_n454_), .A3(new_n1524_), .ZN(new_n1580_));
  NAND3_X1  g1266(.A1(new_n1579_), .A2(new_n1580_), .A3(new_n1452_), .ZN(new_n1581_));
  AOI21_X1  g1267(.A(new_n1575_), .B1(new_n1578_), .B2(new_n1581_), .ZN(new_n1582_));
  NOR2_X1   g1268(.A1(new_n1574_), .A2(new_n1582_), .ZN(G321));
  INV_X1    g1269(.A(new_n1305_), .ZN(new_n1584_));
  NAND4_X1  g1270(.A1(new_n404_), .A2(new_n397_), .A3(new_n388_), .A4(new_n393_), .ZN(new_n1585_));
  NAND4_X1  g1271(.A1(new_n1585_), .A2(new_n1341_), .A3(new_n664_), .A4(new_n1339_), .ZN(new_n1586_));
  NOR2_X1   g1272(.A1(new_n1586_), .A2(new_n656_), .ZN(new_n1587_));
  INV_X1    g1273(.A(new_n395_), .ZN(new_n1588_));
  OAI211_X1 g1274(.A(new_n388_), .B(new_n393_), .C1(new_n396_), .C2(new_n1588_), .ZN(new_n1589_));
  NAND3_X1  g1275(.A1(new_n1589_), .A2(new_n653_), .A3(new_n1346_), .ZN(new_n1590_));
  NOR2_X1   g1276(.A1(new_n1588_), .A2(new_n396_), .ZN(new_n1591_));
  INV_X1    g1277(.A(new_n1591_), .ZN(new_n1592_));
  NAND2_X1  g1278(.A1(new_n1590_), .A2(new_n1592_), .ZN(new_n1593_));
  NOR2_X1   g1279(.A1(new_n1347_), .A2(new_n661_), .ZN(new_n1594_));
  NAND2_X1  g1280(.A1(new_n397_), .A2(new_n393_), .ZN(new_n1595_));
  NAND2_X1  g1281(.A1(new_n1594_), .A2(new_n1595_), .ZN(new_n1596_));
  NAND4_X1  g1282(.A1(new_n1589_), .A2(new_n653_), .A3(new_n1346_), .A4(new_n1591_), .ZN(new_n1597_));
  AND3_X1   g1283(.A1(new_n1593_), .A2(new_n1596_), .A3(new_n1597_), .ZN(new_n1598_));
  AOI21_X1  g1284(.A(new_n1596_), .B1(new_n1593_), .B2(new_n1597_), .ZN(new_n1599_));
  OAI21_X1  g1285(.A(new_n1587_), .B1(new_n1598_), .B2(new_n1599_), .ZN(new_n1600_));
  NAND2_X1  g1286(.A1(new_n1593_), .A2(new_n1597_), .ZN(new_n1601_));
  INV_X1    g1287(.A(new_n1596_), .ZN(new_n1602_));
  NAND2_X1  g1288(.A1(new_n1601_), .A2(new_n1602_), .ZN(new_n1603_));
  OR2_X1    g1289(.A1(new_n1586_), .A2(new_n656_), .ZN(new_n1604_));
  NAND3_X1  g1290(.A1(new_n1593_), .A2(new_n1596_), .A3(new_n1597_), .ZN(new_n1605_));
  NAND3_X1  g1291(.A1(new_n1603_), .A2(new_n1604_), .A3(new_n1605_), .ZN(new_n1606_));
  AND3_X1   g1292(.A1(new_n1600_), .A2(new_n1606_), .A3(new_n397_), .ZN(new_n1607_));
  AOI21_X1  g1293(.A(new_n397_), .B1(new_n1600_), .B2(new_n1606_), .ZN(new_n1608_));
  OAI21_X1  g1294(.A(new_n982_), .B1(new_n1607_), .B2(new_n1608_), .ZN(new_n1609_));
  NOR3_X1   g1295(.A1(new_n1598_), .A2(new_n1599_), .A3(new_n1587_), .ZN(new_n1610_));
  AOI21_X1  g1296(.A(new_n1604_), .B1(new_n1603_), .B2(new_n1605_), .ZN(new_n1611_));
  OAI21_X1  g1297(.A(new_n398_), .B1(new_n1610_), .B2(new_n1611_), .ZN(new_n1612_));
  NAND3_X1  g1298(.A1(new_n1600_), .A2(new_n1606_), .A3(new_n397_), .ZN(new_n1613_));
  NAND3_X1  g1299(.A1(new_n1612_), .A2(new_n393_), .A3(new_n1613_), .ZN(new_n1614_));
  AND3_X1   g1300(.A1(new_n1609_), .A2(new_n382_), .A3(new_n1614_), .ZN(new_n1615_));
  AOI21_X1  g1301(.A(new_n382_), .B1(new_n1609_), .B2(new_n1614_), .ZN(new_n1616_));
  NOR3_X1   g1302(.A1(new_n1615_), .A2(new_n1616_), .A3(new_n1336_), .ZN(new_n1617_));
  NOR3_X1   g1303(.A1(new_n1607_), .A2(new_n1608_), .A3(new_n982_), .ZN(new_n1618_));
  AOI21_X1  g1304(.A(new_n393_), .B1(new_n1612_), .B2(new_n1613_), .ZN(new_n1619_));
  OAI21_X1  g1305(.A(new_n381_), .B1(new_n1618_), .B2(new_n1619_), .ZN(new_n1620_));
  NAND3_X1  g1306(.A1(new_n1609_), .A2(new_n1614_), .A3(new_n382_), .ZN(new_n1621_));
  AOI21_X1  g1307(.A(new_n388_), .B1(new_n1620_), .B2(new_n1621_), .ZN(new_n1622_));
  OAI21_X1  g1308(.A(new_n405_), .B1(new_n1617_), .B2(new_n1622_), .ZN(new_n1623_));
  OAI21_X1  g1309(.A(new_n1336_), .B1(new_n1615_), .B2(new_n1616_), .ZN(new_n1624_));
  NAND3_X1  g1310(.A1(new_n1620_), .A2(new_n388_), .A3(new_n1621_), .ZN(new_n1625_));
  NAND3_X1  g1311(.A1(new_n1624_), .A2(new_n404_), .A3(new_n1625_), .ZN(new_n1626_));
  AOI21_X1  g1312(.A(new_n1584_), .B1(new_n1623_), .B2(new_n1626_), .ZN(new_n1627_));
  NAND4_X1  g1313(.A1(new_n1341_), .A2(new_n1339_), .A3(new_n664_), .A4(new_n655_), .ZN(new_n1628_));
  OAI211_X1 g1314(.A(new_n1346_), .B(new_n653_), .C1(new_n1354_), .C2(new_n1336_), .ZN(new_n1629_));
  NAND2_X1  g1315(.A1(new_n1629_), .A2(new_n1340_), .ZN(new_n1630_));
  AOI21_X1  g1316(.A(new_n654_), .B1(new_n1347_), .B2(new_n388_), .ZN(new_n1631_));
  NAND3_X1  g1317(.A1(new_n1631_), .A2(new_n647_), .A3(new_n1346_), .ZN(new_n1632_));
  AND3_X1   g1318(.A1(new_n1630_), .A2(new_n1632_), .A3(new_n1594_), .ZN(new_n1633_));
  AOI21_X1  g1319(.A(new_n1594_), .B1(new_n1630_), .B2(new_n1632_), .ZN(new_n1634_));
  OAI21_X1  g1320(.A(new_n1628_), .B1(new_n1633_), .B2(new_n1634_), .ZN(new_n1635_));
  NAND2_X1  g1321(.A1(new_n1630_), .A2(new_n1632_), .ZN(new_n1636_));
  NAND2_X1  g1322(.A1(new_n1354_), .A2(new_n660_), .ZN(new_n1637_));
  NAND2_X1  g1323(.A1(new_n1636_), .A2(new_n1637_), .ZN(new_n1638_));
  INV_X1    g1324(.A(new_n1628_), .ZN(new_n1639_));
  NAND3_X1  g1325(.A1(new_n1630_), .A2(new_n1632_), .A3(new_n1594_), .ZN(new_n1640_));
  NAND3_X1  g1326(.A1(new_n1638_), .A2(new_n1639_), .A3(new_n1640_), .ZN(new_n1641_));
  AND3_X1   g1327(.A1(new_n1635_), .A2(new_n1641_), .A3(new_n397_), .ZN(new_n1642_));
  AOI21_X1  g1328(.A(new_n397_), .B1(new_n1635_), .B2(new_n1641_), .ZN(new_n1643_));
  OAI21_X1  g1329(.A(new_n982_), .B1(new_n1642_), .B2(new_n1643_), .ZN(new_n1644_));
  NOR3_X1   g1330(.A1(new_n1633_), .A2(new_n1634_), .A3(new_n1628_), .ZN(new_n1645_));
  AOI21_X1  g1331(.A(new_n1639_), .B1(new_n1638_), .B2(new_n1640_), .ZN(new_n1646_));
  OAI21_X1  g1332(.A(new_n398_), .B1(new_n1645_), .B2(new_n1646_), .ZN(new_n1647_));
  NAND3_X1  g1333(.A1(new_n1635_), .A2(new_n1641_), .A3(new_n397_), .ZN(new_n1648_));
  NAND3_X1  g1334(.A1(new_n1647_), .A2(new_n393_), .A3(new_n1648_), .ZN(new_n1649_));
  AND3_X1   g1335(.A1(new_n1644_), .A2(new_n382_), .A3(new_n1649_), .ZN(new_n1650_));
  AOI21_X1  g1336(.A(new_n382_), .B1(new_n1644_), .B2(new_n1649_), .ZN(new_n1651_));
  OAI21_X1  g1337(.A(new_n1336_), .B1(new_n1650_), .B2(new_n1651_), .ZN(new_n1652_));
  NOR3_X1   g1338(.A1(new_n1642_), .A2(new_n1643_), .A3(new_n982_), .ZN(new_n1653_));
  AOI21_X1  g1339(.A(new_n393_), .B1(new_n1647_), .B2(new_n1648_), .ZN(new_n1654_));
  OAI21_X1  g1340(.A(new_n381_), .B1(new_n1653_), .B2(new_n1654_), .ZN(new_n1655_));
  NAND3_X1  g1341(.A1(new_n1644_), .A2(new_n1649_), .A3(new_n382_), .ZN(new_n1656_));
  NAND3_X1  g1342(.A1(new_n1655_), .A2(new_n388_), .A3(new_n1656_), .ZN(new_n1657_));
  AND3_X1   g1343(.A1(new_n1652_), .A2(new_n404_), .A3(new_n1657_), .ZN(new_n1658_));
  AOI21_X1  g1344(.A(new_n404_), .B1(new_n1652_), .B2(new_n1657_), .ZN(new_n1659_));
  NOR3_X1   g1345(.A1(new_n1658_), .A2(new_n1659_), .A3(new_n1305_), .ZN(new_n1660_));
  NAND2_X1  g1346(.A1(new_n407_), .A2(G38), .ZN(new_n1661_));
  XOR2_X1   g1347(.A(new_n410_), .B(new_n1661_), .Z(new_n1662_));
  INV_X1    g1348(.A(new_n1662_), .ZN(new_n1663_));
  NAND3_X1  g1349(.A1(new_n1584_), .A2(new_n667_), .A3(new_n1663_), .ZN(new_n1664_));
  NOR2_X1   g1350(.A1(new_n407_), .A2(G38), .ZN(new_n1665_));
  XNOR2_X1  g1351(.A(new_n410_), .B(new_n1665_), .ZN(new_n1666_));
  INV_X1    g1352(.A(new_n1666_), .ZN(new_n1667_));
  NAND3_X1  g1353(.A1(new_n1584_), .A2(new_n666_), .A3(new_n1667_), .ZN(new_n1668_));
  OAI211_X1 g1354(.A(new_n1305_), .B(new_n1663_), .C1(new_n667_), .C2(new_n983_), .ZN(new_n1669_));
  NAND4_X1  g1355(.A1(new_n1305_), .A2(new_n666_), .A3(new_n984_), .A4(new_n1667_), .ZN(new_n1670_));
  NAND4_X1  g1356(.A1(new_n1664_), .A2(new_n1668_), .A3(new_n1669_), .A4(new_n1670_), .ZN(new_n1671_));
  INV_X1    g1357(.A(new_n1671_), .ZN(new_n1672_));
  NOR3_X1   g1358(.A1(new_n1627_), .A2(new_n1660_), .A3(new_n1672_), .ZN(new_n1673_));
  AND3_X1   g1359(.A1(new_n1624_), .A2(new_n404_), .A3(new_n1625_), .ZN(new_n1674_));
  AOI21_X1  g1360(.A(new_n404_), .B1(new_n1624_), .B2(new_n1625_), .ZN(new_n1675_));
  OAI21_X1  g1361(.A(new_n1305_), .B1(new_n1674_), .B2(new_n1675_), .ZN(new_n1676_));
  INV_X1    g1362(.A(new_n1659_), .ZN(new_n1677_));
  NAND3_X1  g1363(.A1(new_n1652_), .A2(new_n404_), .A3(new_n1657_), .ZN(new_n1678_));
  NAND3_X1  g1364(.A1(new_n1677_), .A2(new_n1584_), .A3(new_n1678_), .ZN(new_n1679_));
  AOI21_X1  g1365(.A(new_n1671_), .B1(new_n1676_), .B2(new_n1679_), .ZN(new_n1680_));
  NOR2_X1   g1366(.A1(new_n1673_), .A2(new_n1680_), .ZN(G338));
  AOI21_X1  g1367(.A(new_n507_), .B1(G4526), .B2(new_n996_), .ZN(new_n1682_));
  OAI21_X1  g1368(.A(new_n548_), .B1(new_n1682_), .B2(new_n968_), .ZN(new_n1683_));
  INV_X1    g1369(.A(new_n1683_), .ZN(new_n1684_));
  NAND4_X1  g1370(.A1(new_n604_), .A2(new_n585_), .A3(new_n592_), .A4(new_n599_), .ZN(new_n1685_));
  NAND4_X1  g1371(.A1(new_n1685_), .A2(new_n1407_), .A3(new_n684_), .A4(new_n1406_), .ZN(new_n1686_));
  NOR2_X1   g1372(.A1(new_n1686_), .A2(new_n677_), .ZN(new_n1687_));
  INV_X1    g1373(.A(G4394), .ZN(new_n1688_));
  OAI211_X1 g1374(.A(new_n592_), .B(new_n599_), .C1(new_n1688_), .C2(new_n603_), .ZN(new_n1689_));
  NAND3_X1  g1375(.A1(new_n1689_), .A2(new_n1412_), .A3(new_n1413_), .ZN(new_n1690_));
  INV_X1    g1376(.A(new_n603_), .ZN(new_n1691_));
  NAND2_X1  g1377(.A1(new_n1691_), .A2(G4394), .ZN(new_n1692_));
  NAND2_X1  g1378(.A1(new_n1690_), .A2(new_n1692_), .ZN(new_n1693_));
  NAND2_X1  g1379(.A1(new_n1421_), .A2(new_n1418_), .ZN(new_n1694_));
  INV_X1    g1380(.A(new_n1694_), .ZN(new_n1695_));
  OAI21_X1  g1381(.A(new_n1695_), .B1(new_n1403_), .B2(new_n605_), .ZN(new_n1696_));
  INV_X1    g1382(.A(new_n1692_), .ZN(new_n1697_));
  NAND4_X1  g1383(.A1(new_n1689_), .A2(new_n1412_), .A3(new_n1413_), .A4(new_n1697_), .ZN(new_n1698_));
  AND3_X1   g1384(.A1(new_n1693_), .A2(new_n1696_), .A3(new_n1698_), .ZN(new_n1699_));
  AOI21_X1  g1385(.A(new_n1696_), .B1(new_n1693_), .B2(new_n1698_), .ZN(new_n1700_));
  OAI21_X1  g1386(.A(new_n1687_), .B1(new_n1699_), .B2(new_n1700_), .ZN(new_n1701_));
  NAND2_X1  g1387(.A1(new_n1693_), .A2(new_n1698_), .ZN(new_n1702_));
  INV_X1    g1388(.A(new_n1696_), .ZN(new_n1703_));
  NAND2_X1  g1389(.A1(new_n1702_), .A2(new_n1703_), .ZN(new_n1704_));
  OR2_X1    g1390(.A1(new_n1686_), .A2(new_n677_), .ZN(new_n1705_));
  NAND3_X1  g1391(.A1(new_n1693_), .A2(new_n1696_), .A3(new_n1698_), .ZN(new_n1706_));
  NAND3_X1  g1392(.A1(new_n1704_), .A2(new_n1705_), .A3(new_n1706_), .ZN(new_n1707_));
  AND3_X1   g1393(.A1(new_n1701_), .A2(new_n1707_), .A3(new_n604_), .ZN(new_n1708_));
  AOI21_X1  g1394(.A(new_n604_), .B1(new_n1701_), .B2(new_n1707_), .ZN(new_n1709_));
  OAI21_X1  g1395(.A(new_n1403_), .B1(new_n1708_), .B2(new_n1709_), .ZN(new_n1710_));
  NOR3_X1   g1396(.A1(new_n1699_), .A2(new_n1700_), .A3(new_n1687_), .ZN(new_n1711_));
  AOI21_X1  g1397(.A(new_n1705_), .B1(new_n1704_), .B2(new_n1706_), .ZN(new_n1712_));
  OAI21_X1  g1398(.A(new_n605_), .B1(new_n1711_), .B2(new_n1712_), .ZN(new_n1713_));
  NAND3_X1  g1399(.A1(new_n1701_), .A2(new_n1707_), .A3(new_n604_), .ZN(new_n1714_));
  NAND3_X1  g1400(.A1(new_n1713_), .A2(new_n599_), .A3(new_n1714_), .ZN(new_n1715_));
  AND3_X1   g1401(.A1(new_n1710_), .A2(new_n578_), .A3(new_n1715_), .ZN(new_n1716_));
  AOI21_X1  g1402(.A(new_n578_), .B1(new_n1710_), .B2(new_n1715_), .ZN(new_n1717_));
  NOR3_X1   g1403(.A1(new_n1716_), .A2(new_n1717_), .A3(new_n973_), .ZN(new_n1718_));
  NOR3_X1   g1404(.A1(new_n1708_), .A2(new_n1709_), .A3(new_n1403_), .ZN(new_n1719_));
  AOI21_X1  g1405(.A(new_n599_), .B1(new_n1713_), .B2(new_n1714_), .ZN(new_n1720_));
  OAI21_X1  g1406(.A(new_n683_), .B1(new_n1719_), .B2(new_n1720_), .ZN(new_n1721_));
  NAND3_X1  g1407(.A1(new_n1710_), .A2(new_n1715_), .A3(new_n578_), .ZN(new_n1722_));
  AOI21_X1  g1408(.A(new_n592_), .B1(new_n1721_), .B2(new_n1722_), .ZN(new_n1723_));
  OAI21_X1  g1409(.A(new_n669_), .B1(new_n1718_), .B2(new_n1723_), .ZN(new_n1724_));
  OAI21_X1  g1410(.A(new_n973_), .B1(new_n1716_), .B2(new_n1717_), .ZN(new_n1725_));
  NAND3_X1  g1411(.A1(new_n1721_), .A2(new_n592_), .A3(new_n1722_), .ZN(new_n1726_));
  NAND3_X1  g1412(.A1(new_n1725_), .A2(new_n585_), .A3(new_n1726_), .ZN(new_n1727_));
  AOI21_X1  g1413(.A(new_n1684_), .B1(new_n1724_), .B2(new_n1727_), .ZN(new_n1728_));
  NAND4_X1  g1414(.A1(new_n1407_), .A2(new_n676_), .A3(new_n1406_), .A4(new_n684_), .ZN(new_n1729_));
  OAI211_X1 g1415(.A(new_n1412_), .B(new_n1413_), .C1(new_n1421_), .C2(new_n973_), .ZN(new_n1730_));
  NAND2_X1  g1416(.A1(new_n1730_), .A2(new_n670_), .ZN(new_n1731_));
  NAND4_X1  g1417(.A1(new_n1414_), .A2(new_n1412_), .A3(new_n671_), .A4(new_n1413_), .ZN(new_n1732_));
  AND3_X1   g1418(.A1(new_n1731_), .A2(new_n1695_), .A3(new_n1732_), .ZN(new_n1733_));
  AOI21_X1  g1419(.A(new_n1695_), .B1(new_n1731_), .B2(new_n1732_), .ZN(new_n1734_));
  OAI21_X1  g1420(.A(new_n1729_), .B1(new_n1733_), .B2(new_n1734_), .ZN(new_n1735_));
  NAND2_X1  g1421(.A1(new_n1731_), .A2(new_n1732_), .ZN(new_n1736_));
  NAND2_X1  g1422(.A1(new_n1736_), .A2(new_n1694_), .ZN(new_n1737_));
  INV_X1    g1423(.A(new_n1729_), .ZN(new_n1738_));
  NAND3_X1  g1424(.A1(new_n1731_), .A2(new_n1695_), .A3(new_n1732_), .ZN(new_n1739_));
  NAND3_X1  g1425(.A1(new_n1737_), .A2(new_n1738_), .A3(new_n1739_), .ZN(new_n1740_));
  AND3_X1   g1426(.A1(new_n1735_), .A2(new_n1740_), .A3(new_n604_), .ZN(new_n1741_));
  AOI21_X1  g1427(.A(new_n604_), .B1(new_n1735_), .B2(new_n1740_), .ZN(new_n1742_));
  OAI21_X1  g1428(.A(new_n1403_), .B1(new_n1741_), .B2(new_n1742_), .ZN(new_n1743_));
  NOR3_X1   g1429(.A1(new_n1733_), .A2(new_n1734_), .A3(new_n1729_), .ZN(new_n1744_));
  AOI21_X1  g1430(.A(new_n1738_), .B1(new_n1737_), .B2(new_n1739_), .ZN(new_n1745_));
  OAI21_X1  g1431(.A(new_n605_), .B1(new_n1744_), .B2(new_n1745_), .ZN(new_n1746_));
  NAND3_X1  g1432(.A1(new_n1735_), .A2(new_n1740_), .A3(new_n604_), .ZN(new_n1747_));
  NAND3_X1  g1433(.A1(new_n1746_), .A2(new_n599_), .A3(new_n1747_), .ZN(new_n1748_));
  AND3_X1   g1434(.A1(new_n1743_), .A2(new_n578_), .A3(new_n1748_), .ZN(new_n1749_));
  AOI21_X1  g1435(.A(new_n578_), .B1(new_n1743_), .B2(new_n1748_), .ZN(new_n1750_));
  OAI21_X1  g1436(.A(new_n973_), .B1(new_n1749_), .B2(new_n1750_), .ZN(new_n1751_));
  NOR3_X1   g1437(.A1(new_n1741_), .A2(new_n1742_), .A3(new_n1403_), .ZN(new_n1752_));
  AOI21_X1  g1438(.A(new_n599_), .B1(new_n1746_), .B2(new_n1747_), .ZN(new_n1753_));
  OAI21_X1  g1439(.A(new_n683_), .B1(new_n1752_), .B2(new_n1753_), .ZN(new_n1754_));
  NAND3_X1  g1440(.A1(new_n1743_), .A2(new_n1748_), .A3(new_n578_), .ZN(new_n1755_));
  NAND3_X1  g1441(.A1(new_n1754_), .A2(new_n592_), .A3(new_n1755_), .ZN(new_n1756_));
  AND3_X1   g1442(.A1(new_n1751_), .A2(new_n585_), .A3(new_n1756_), .ZN(new_n1757_));
  AOI21_X1  g1443(.A(new_n585_), .B1(new_n1751_), .B2(new_n1756_), .ZN(new_n1758_));
  NOR3_X1   g1444(.A1(new_n1757_), .A2(new_n1758_), .A3(new_n1683_), .ZN(new_n1759_));
  OAI22_X1  g1445(.A1(new_n571_), .A2(new_n572_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n1760_));
  OAI211_X1 g1446(.A(new_n691_), .B(G4420), .C1(G4427), .C2(new_n558_), .ZN(new_n1761_));
  NAND3_X1  g1447(.A1(new_n1431_), .A2(new_n1760_), .A3(new_n1761_), .ZN(new_n1762_));
  NAND2_X1  g1448(.A1(new_n1761_), .A2(new_n1760_), .ZN(new_n1763_));
  NAND4_X1  g1449(.A1(new_n1430_), .A2(new_n689_), .A3(new_n695_), .A4(new_n1763_), .ZN(new_n1764_));
  AOI21_X1  g1450(.A(new_n977_), .B1(new_n1762_), .B2(new_n1764_), .ZN(new_n1765_));
  INV_X1    g1451(.A(new_n1765_), .ZN(new_n1766_));
  NAND3_X1  g1452(.A1(new_n1762_), .A2(new_n977_), .A3(new_n1764_), .ZN(new_n1767_));
  AOI21_X1  g1453(.A(new_n562_), .B1(new_n1766_), .B2(new_n1767_), .ZN(new_n1768_));
  INV_X1    g1454(.A(new_n1767_), .ZN(new_n1769_));
  NOR3_X1   g1455(.A1(new_n1769_), .A2(new_n1765_), .A3(new_n563_), .ZN(new_n1770_));
  OAI21_X1  g1456(.A(new_n568_), .B1(new_n1768_), .B2(new_n1770_), .ZN(new_n1771_));
  OAI21_X1  g1457(.A(new_n563_), .B1(new_n1769_), .B2(new_n1765_), .ZN(new_n1772_));
  NAND3_X1  g1458(.A1(new_n1766_), .A2(new_n562_), .A3(new_n1767_), .ZN(new_n1773_));
  NAND3_X1  g1459(.A1(new_n1772_), .A2(new_n1773_), .A3(new_n976_), .ZN(new_n1774_));
  AND3_X1   g1460(.A1(new_n1771_), .A2(new_n553_), .A3(new_n1774_), .ZN(new_n1775_));
  AOI21_X1  g1461(.A(new_n553_), .B1(new_n1771_), .B2(new_n1774_), .ZN(new_n1776_));
  OAI211_X1 g1462(.A(new_n686_), .B(new_n1684_), .C1(new_n1775_), .C2(new_n1776_), .ZN(new_n1777_));
  INV_X1    g1463(.A(new_n686_), .ZN(new_n1778_));
  NAND3_X1  g1464(.A1(new_n553_), .A2(new_n562_), .A3(new_n692_), .ZN(new_n1779_));
  NAND3_X1  g1465(.A1(new_n1779_), .A2(new_n689_), .A3(new_n695_), .ZN(new_n1780_));
  OAI21_X1  g1466(.A(new_n1442_), .B1(new_n558_), .B2(G4427), .ZN(new_n1781_));
  OAI21_X1  g1467(.A(new_n692_), .B1(new_n559_), .B2(new_n557_), .ZN(new_n1782_));
  NAND2_X1  g1468(.A1(new_n1781_), .A2(new_n1782_), .ZN(new_n1783_));
  OR2_X1    g1469(.A1(new_n1780_), .A2(new_n1783_), .ZN(new_n1784_));
  NAND2_X1  g1470(.A1(new_n1780_), .A2(new_n1783_), .ZN(new_n1785_));
  NAND3_X1  g1471(.A1(new_n1784_), .A2(new_n977_), .A3(new_n1785_), .ZN(new_n1786_));
  INV_X1    g1472(.A(new_n1786_), .ZN(new_n1787_));
  AOI21_X1  g1473(.A(new_n977_), .B1(new_n1784_), .B2(new_n1785_), .ZN(new_n1788_));
  NOR3_X1   g1474(.A1(new_n1787_), .A2(new_n1788_), .A3(new_n563_), .ZN(new_n1789_));
  NAND2_X1  g1475(.A1(new_n1784_), .A2(new_n1785_), .ZN(new_n1790_));
  NAND2_X1  g1476(.A1(new_n1790_), .A2(new_n573_), .ZN(new_n1791_));
  AOI21_X1  g1477(.A(new_n562_), .B1(new_n1791_), .B2(new_n1786_), .ZN(new_n1792_));
  OAI21_X1  g1478(.A(new_n568_), .B1(new_n1789_), .B2(new_n1792_), .ZN(new_n1793_));
  OAI21_X1  g1479(.A(new_n563_), .B1(new_n1787_), .B2(new_n1788_), .ZN(new_n1794_));
  NAND3_X1  g1480(.A1(new_n1791_), .A2(new_n1786_), .A3(new_n562_), .ZN(new_n1795_));
  NAND3_X1  g1481(.A1(new_n1794_), .A2(new_n976_), .A3(new_n1795_), .ZN(new_n1796_));
  AND3_X1   g1482(.A1(new_n1793_), .A2(new_n553_), .A3(new_n1796_), .ZN(new_n1797_));
  AOI21_X1  g1483(.A(new_n553_), .B1(new_n1793_), .B2(new_n1796_), .ZN(new_n1798_));
  OAI211_X1 g1484(.A(new_n1778_), .B(new_n1684_), .C1(new_n1797_), .C2(new_n1798_), .ZN(new_n1799_));
  NAND2_X1  g1485(.A1(new_n1778_), .A2(new_n975_), .ZN(new_n1800_));
  INV_X1    g1486(.A(new_n1800_), .ZN(new_n1801_));
  OAI211_X1 g1487(.A(new_n1683_), .B(new_n1801_), .C1(new_n1797_), .C2(new_n1798_), .ZN(new_n1802_));
  OAI211_X1 g1488(.A(new_n1683_), .B(new_n1800_), .C1(new_n1775_), .C2(new_n1776_), .ZN(new_n1803_));
  AND4_X1   g1489(.A1(new_n1777_), .A2(new_n1799_), .A3(new_n1802_), .A4(new_n1803_), .ZN(new_n1804_));
  NOR3_X1   g1490(.A1(new_n1728_), .A2(new_n1759_), .A3(new_n1804_), .ZN(new_n1805_));
  NAND4_X1  g1491(.A1(new_n1777_), .A2(new_n1799_), .A3(new_n1802_), .A4(new_n1803_), .ZN(new_n1806_));
  AND3_X1   g1492(.A1(new_n1725_), .A2(new_n585_), .A3(new_n1726_), .ZN(new_n1807_));
  AOI21_X1  g1493(.A(new_n585_), .B1(new_n1725_), .B2(new_n1726_), .ZN(new_n1808_));
  OAI21_X1  g1494(.A(new_n1683_), .B1(new_n1807_), .B2(new_n1808_), .ZN(new_n1809_));
  INV_X1    g1495(.A(new_n1758_), .ZN(new_n1810_));
  NAND3_X1  g1496(.A1(new_n1751_), .A2(new_n585_), .A3(new_n1756_), .ZN(new_n1811_));
  NAND3_X1  g1497(.A1(new_n1810_), .A2(new_n1811_), .A3(new_n1684_), .ZN(new_n1812_));
  AOI21_X1  g1498(.A(new_n1806_), .B1(new_n1809_), .B2(new_n1812_), .ZN(new_n1813_));
  NOR2_X1   g1499(.A1(new_n1805_), .A2(new_n1813_), .ZN(G370));
  NAND4_X1  g1500(.A1(new_n470_), .A2(new_n374_), .A3(new_n481_), .A4(new_n488_), .ZN(new_n1815_));
  NAND4_X1  g1501(.A1(new_n1815_), .A2(new_n1010_), .A3(new_n504_), .A4(new_n1008_), .ZN(new_n1816_));
  NOR2_X1   g1502(.A1(new_n1816_), .A2(new_n498_), .ZN(new_n1817_));
  OAI211_X1 g1503(.A(new_n481_), .B(new_n488_), .C1(new_n472_), .C2(new_n373_), .ZN(new_n1818_));
  NAND3_X1  g1504(.A1(new_n1818_), .A2(new_n1019_), .A3(new_n1022_), .ZN(new_n1819_));
  NOR2_X1   g1505(.A1(new_n472_), .A2(new_n373_), .ZN(new_n1820_));
  INV_X1    g1506(.A(new_n1820_), .ZN(new_n1821_));
  NAND2_X1  g1507(.A1(new_n1819_), .A2(new_n1821_), .ZN(new_n1822_));
  NOR2_X1   g1508(.A1(new_n1016_), .A2(new_n501_), .ZN(new_n1823_));
  OAI21_X1  g1509(.A(new_n1823_), .B1(new_n611_), .B2(new_n995_), .ZN(new_n1824_));
  NAND4_X1  g1510(.A1(new_n1818_), .A2(new_n1019_), .A3(new_n1022_), .A4(new_n1820_), .ZN(new_n1825_));
  AND3_X1   g1511(.A1(new_n1822_), .A2(new_n1824_), .A3(new_n1825_), .ZN(new_n1826_));
  AOI21_X1  g1512(.A(new_n1824_), .B1(new_n1822_), .B2(new_n1825_), .ZN(new_n1827_));
  OAI21_X1  g1513(.A(new_n1817_), .B1(new_n1826_), .B2(new_n1827_), .ZN(new_n1828_));
  NAND2_X1  g1514(.A1(new_n1822_), .A2(new_n1825_), .ZN(new_n1829_));
  INV_X1    g1515(.A(new_n1824_), .ZN(new_n1830_));
  NAND2_X1  g1516(.A1(new_n1829_), .A2(new_n1830_), .ZN(new_n1831_));
  OR2_X1    g1517(.A1(new_n1816_), .A2(new_n498_), .ZN(new_n1832_));
  NAND3_X1  g1518(.A1(new_n1822_), .A2(new_n1824_), .A3(new_n1825_), .ZN(new_n1833_));
  NAND3_X1  g1519(.A1(new_n1831_), .A2(new_n1832_), .A3(new_n1833_), .ZN(new_n1834_));
  AND3_X1   g1520(.A1(new_n1828_), .A2(new_n1834_), .A3(new_n374_), .ZN(new_n1835_));
  AOI21_X1  g1521(.A(new_n374_), .B1(new_n1828_), .B2(new_n1834_), .ZN(new_n1836_));
  OAI21_X1  g1522(.A(new_n995_), .B1(new_n1835_), .B2(new_n1836_), .ZN(new_n1837_));
  NOR3_X1   g1523(.A1(new_n1826_), .A2(new_n1827_), .A3(new_n1817_), .ZN(new_n1838_));
  AOI21_X1  g1524(.A(new_n1832_), .B1(new_n1831_), .B2(new_n1833_), .ZN(new_n1839_));
  OAI21_X1  g1525(.A(new_n611_), .B1(new_n1838_), .B2(new_n1839_), .ZN(new_n1840_));
  NAND3_X1  g1526(.A1(new_n1828_), .A2(new_n1834_), .A3(new_n374_), .ZN(new_n1841_));
  NAND3_X1  g1527(.A1(new_n1840_), .A2(new_n488_), .A3(new_n1841_), .ZN(new_n1842_));
  AND3_X1   g1528(.A1(new_n1837_), .A2(new_n494_), .A3(new_n1842_), .ZN(new_n1843_));
  AOI21_X1  g1529(.A(new_n494_), .B1(new_n1837_), .B2(new_n1842_), .ZN(new_n1844_));
  NOR3_X1   g1530(.A1(new_n1843_), .A2(new_n1844_), .A3(new_n1031_), .ZN(new_n1845_));
  NOR3_X1   g1531(.A1(new_n1835_), .A2(new_n1836_), .A3(new_n995_), .ZN(new_n1846_));
  AOI21_X1  g1532(.A(new_n488_), .B1(new_n1840_), .B2(new_n1841_), .ZN(new_n1847_));
  OAI21_X1  g1533(.A(new_n493_), .B1(new_n1846_), .B2(new_n1847_), .ZN(new_n1848_));
  NAND3_X1  g1534(.A1(new_n1837_), .A2(new_n1842_), .A3(new_n494_), .ZN(new_n1849_));
  AOI21_X1  g1535(.A(new_n481_), .B1(new_n1848_), .B2(new_n1849_), .ZN(new_n1850_));
  OAI21_X1  g1536(.A(new_n471_), .B1(new_n1845_), .B2(new_n1850_), .ZN(new_n1851_));
  OAI21_X1  g1537(.A(new_n1031_), .B1(new_n1843_), .B2(new_n1844_), .ZN(new_n1852_));
  NAND3_X1  g1538(.A1(new_n1848_), .A2(new_n481_), .A3(new_n1849_), .ZN(new_n1853_));
  NAND3_X1  g1539(.A1(new_n1852_), .A2(new_n470_), .A3(new_n1853_), .ZN(new_n1854_));
  AOI21_X1  g1540(.A(new_n375_), .B1(new_n1851_), .B2(new_n1854_), .ZN(new_n1855_));
  NAND4_X1  g1541(.A1(new_n1010_), .A2(new_n497_), .A3(new_n1008_), .A4(new_n504_), .ZN(new_n1856_));
  OAI211_X1 g1542(.A(new_n1019_), .B(new_n1022_), .C1(new_n1029_), .C2(new_n1031_), .ZN(new_n1857_));
  NAND2_X1  g1543(.A1(new_n1857_), .A2(new_n1009_), .ZN(new_n1858_));
  NAND4_X1  g1544(.A1(new_n1017_), .A2(new_n1019_), .A3(new_n473_), .A4(new_n1022_), .ZN(new_n1859_));
  AND3_X1   g1545(.A1(new_n1858_), .A2(new_n1859_), .A3(new_n1823_), .ZN(new_n1860_));
  AOI21_X1  g1546(.A(new_n1823_), .B1(new_n1858_), .B2(new_n1859_), .ZN(new_n1861_));
  OAI21_X1  g1547(.A(new_n1856_), .B1(new_n1860_), .B2(new_n1861_), .ZN(new_n1862_));
  NAND2_X1  g1548(.A1(new_n1858_), .A2(new_n1859_), .ZN(new_n1863_));
  INV_X1    g1549(.A(new_n1823_), .ZN(new_n1864_));
  NAND2_X1  g1550(.A1(new_n1863_), .A2(new_n1864_), .ZN(new_n1865_));
  INV_X1    g1551(.A(new_n1856_), .ZN(new_n1866_));
  NAND3_X1  g1552(.A1(new_n1858_), .A2(new_n1859_), .A3(new_n1823_), .ZN(new_n1867_));
  NAND3_X1  g1553(.A1(new_n1865_), .A2(new_n1866_), .A3(new_n1867_), .ZN(new_n1868_));
  AND3_X1   g1554(.A1(new_n1862_), .A2(new_n1868_), .A3(new_n374_), .ZN(new_n1869_));
  AOI21_X1  g1555(.A(new_n374_), .B1(new_n1862_), .B2(new_n1868_), .ZN(new_n1870_));
  OAI21_X1  g1556(.A(new_n995_), .B1(new_n1869_), .B2(new_n1870_), .ZN(new_n1871_));
  NOR3_X1   g1557(.A1(new_n1860_), .A2(new_n1861_), .A3(new_n1856_), .ZN(new_n1872_));
  AOI21_X1  g1558(.A(new_n1866_), .B1(new_n1865_), .B2(new_n1867_), .ZN(new_n1873_));
  OAI21_X1  g1559(.A(new_n611_), .B1(new_n1872_), .B2(new_n1873_), .ZN(new_n1874_));
  NAND3_X1  g1560(.A1(new_n1862_), .A2(new_n1868_), .A3(new_n374_), .ZN(new_n1875_));
  NAND3_X1  g1561(.A1(new_n1874_), .A2(new_n488_), .A3(new_n1875_), .ZN(new_n1876_));
  AND3_X1   g1562(.A1(new_n1871_), .A2(new_n494_), .A3(new_n1876_), .ZN(new_n1877_));
  AOI21_X1  g1563(.A(new_n494_), .B1(new_n1871_), .B2(new_n1876_), .ZN(new_n1878_));
  OAI21_X1  g1564(.A(new_n1031_), .B1(new_n1877_), .B2(new_n1878_), .ZN(new_n1879_));
  NOR3_X1   g1565(.A1(new_n1869_), .A2(new_n1870_), .A3(new_n995_), .ZN(new_n1880_));
  AOI21_X1  g1566(.A(new_n488_), .B1(new_n1874_), .B2(new_n1875_), .ZN(new_n1881_));
  OAI21_X1  g1567(.A(new_n493_), .B1(new_n1880_), .B2(new_n1881_), .ZN(new_n1882_));
  NAND3_X1  g1568(.A1(new_n1871_), .A2(new_n1876_), .A3(new_n494_), .ZN(new_n1883_));
  NAND3_X1  g1569(.A1(new_n1882_), .A2(new_n481_), .A3(new_n1883_), .ZN(new_n1884_));
  AND3_X1   g1570(.A1(new_n1879_), .A2(new_n470_), .A3(new_n1884_), .ZN(new_n1885_));
  AOI21_X1  g1571(.A(new_n470_), .B1(new_n1879_), .B2(new_n1884_), .ZN(new_n1886_));
  NOR3_X1   g1572(.A1(new_n1885_), .A2(new_n1886_), .A3(G4526), .ZN(new_n1887_));
  OAI22_X1  g1573(.A1(new_n524_), .A2(new_n525_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n1888_));
  OAI211_X1 g1574(.A(new_n535_), .B(G3729), .C1(G3737), .C2(new_n516_), .ZN(new_n1889_));
  NAND3_X1  g1575(.A1(new_n1041_), .A2(new_n1888_), .A3(new_n1889_), .ZN(new_n1890_));
  NAND2_X1  g1576(.A1(new_n1889_), .A2(new_n1888_), .ZN(new_n1891_));
  NAND4_X1  g1577(.A1(new_n1040_), .A2(new_n544_), .A3(new_n540_), .A4(new_n1891_), .ZN(new_n1892_));
  AOI21_X1  g1578(.A(new_n967_), .B1(new_n1890_), .B2(new_n1892_), .ZN(new_n1893_));
  INV_X1    g1579(.A(new_n1893_), .ZN(new_n1894_));
  NAND3_X1  g1580(.A1(new_n1890_), .A2(new_n967_), .A3(new_n1892_), .ZN(new_n1895_));
  AOI21_X1  g1581(.A(new_n520_), .B1(new_n1894_), .B2(new_n1895_), .ZN(new_n1896_));
  INV_X1    g1582(.A(new_n1895_), .ZN(new_n1897_));
  NOR3_X1   g1583(.A1(new_n1897_), .A2(new_n1893_), .A3(new_n521_), .ZN(new_n1898_));
  OAI21_X1  g1584(.A(new_n531_), .B1(new_n1896_), .B2(new_n1898_), .ZN(new_n1899_));
  OAI21_X1  g1585(.A(new_n521_), .B1(new_n1897_), .B2(new_n1893_), .ZN(new_n1900_));
  NAND3_X1  g1586(.A1(new_n1894_), .A2(new_n520_), .A3(new_n1895_), .ZN(new_n1901_));
  NAND3_X1  g1587(.A1(new_n1900_), .A2(new_n1901_), .A3(new_n534_), .ZN(new_n1902_));
  AND3_X1   g1588(.A1(new_n1899_), .A2(new_n511_), .A3(new_n1902_), .ZN(new_n1903_));
  AOI21_X1  g1589(.A(new_n511_), .B1(new_n1899_), .B2(new_n1902_), .ZN(new_n1904_));
  OAI211_X1 g1590(.A(new_n375_), .B(new_n507_), .C1(new_n1903_), .C2(new_n1904_), .ZN(new_n1905_));
  NAND3_X1  g1591(.A1(new_n511_), .A2(new_n520_), .A3(new_n536_), .ZN(new_n1906_));
  NAND3_X1  g1592(.A1(new_n1906_), .A2(new_n544_), .A3(new_n540_), .ZN(new_n1907_));
  OAI21_X1  g1593(.A(new_n537_), .B1(new_n516_), .B2(G3737), .ZN(new_n1908_));
  OAI21_X1  g1594(.A(new_n536_), .B1(new_n517_), .B2(new_n515_), .ZN(new_n1909_));
  NAND2_X1  g1595(.A1(new_n1908_), .A2(new_n1909_), .ZN(new_n1910_));
  OR2_X1    g1596(.A1(new_n1907_), .A2(new_n1910_), .ZN(new_n1911_));
  NAND2_X1  g1597(.A1(new_n1907_), .A2(new_n1910_), .ZN(new_n1912_));
  NAND3_X1  g1598(.A1(new_n1911_), .A2(new_n967_), .A3(new_n1912_), .ZN(new_n1913_));
  INV_X1    g1599(.A(new_n1913_), .ZN(new_n1914_));
  AOI21_X1  g1600(.A(new_n967_), .B1(new_n1911_), .B2(new_n1912_), .ZN(new_n1915_));
  NOR3_X1   g1601(.A1(new_n1914_), .A2(new_n1915_), .A3(new_n521_), .ZN(new_n1916_));
  NAND2_X1  g1602(.A1(new_n1911_), .A2(new_n1912_), .ZN(new_n1917_));
  NAND2_X1  g1603(.A1(new_n1917_), .A2(new_n526_), .ZN(new_n1918_));
  AOI21_X1  g1604(.A(new_n520_), .B1(new_n1918_), .B2(new_n1913_), .ZN(new_n1919_));
  OAI21_X1  g1605(.A(new_n531_), .B1(new_n1916_), .B2(new_n1919_), .ZN(new_n1920_));
  OAI21_X1  g1606(.A(new_n521_), .B1(new_n1914_), .B2(new_n1915_), .ZN(new_n1921_));
  NAND3_X1  g1607(.A1(new_n1918_), .A2(new_n1913_), .A3(new_n520_), .ZN(new_n1922_));
  NAND3_X1  g1608(.A1(new_n1921_), .A2(new_n534_), .A3(new_n1922_), .ZN(new_n1923_));
  AND3_X1   g1609(.A1(new_n1920_), .A2(new_n511_), .A3(new_n1923_), .ZN(new_n1924_));
  AOI21_X1  g1610(.A(new_n511_), .B1(new_n1920_), .B2(new_n1923_), .ZN(new_n1925_));
  OAI211_X1 g1611(.A(new_n375_), .B(new_n506_), .C1(new_n1924_), .C2(new_n1925_), .ZN(new_n1926_));
  NOR2_X1   g1612(.A1(new_n507_), .A2(new_n996_), .ZN(new_n1927_));
  OAI211_X1 g1613(.A(G4526), .B(new_n1927_), .C1(new_n1924_), .C2(new_n1925_), .ZN(new_n1928_));
  INV_X1    g1614(.A(new_n1927_), .ZN(new_n1929_));
  OAI211_X1 g1615(.A(G4526), .B(new_n1929_), .C1(new_n1903_), .C2(new_n1904_), .ZN(new_n1930_));
  AND4_X1   g1616(.A1(new_n1905_), .A2(new_n1926_), .A3(new_n1928_), .A4(new_n1930_), .ZN(new_n1931_));
  NOR3_X1   g1617(.A1(new_n1855_), .A2(new_n1887_), .A3(new_n1931_), .ZN(new_n1932_));
  NAND4_X1  g1618(.A1(new_n1905_), .A2(new_n1926_), .A3(new_n1928_), .A4(new_n1930_), .ZN(new_n1933_));
  AND3_X1   g1619(.A1(new_n1852_), .A2(new_n470_), .A3(new_n1853_), .ZN(new_n1934_));
  AOI21_X1  g1620(.A(new_n470_), .B1(new_n1852_), .B2(new_n1853_), .ZN(new_n1935_));
  OAI21_X1  g1621(.A(G4526), .B1(new_n1934_), .B2(new_n1935_), .ZN(new_n1936_));
  INV_X1    g1622(.A(new_n1886_), .ZN(new_n1937_));
  NAND3_X1  g1623(.A1(new_n1879_), .A2(new_n470_), .A3(new_n1884_), .ZN(new_n1938_));
  NAND3_X1  g1624(.A1(new_n1937_), .A2(new_n375_), .A3(new_n1938_), .ZN(new_n1939_));
  AOI21_X1  g1625(.A(new_n1933_), .B1(new_n1936_), .B2(new_n1939_), .ZN(new_n1940_));
  NOR2_X1   g1626(.A1(new_n1932_), .A2(new_n1940_), .ZN(G399));
endmodule


