//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_;
  AND2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204_));
  NOR3_X1   g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n202_), .A2(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT10), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT10), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(G99gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  AOI211_X1 g019(.A(new_n220_), .B(G106gat), .C1(new_n214_), .C2(new_n216_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n211_), .B(new_n212_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n226_), .A2(new_n208_), .A3(new_n209_), .A4(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n202_), .A2(new_n203_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n232_), .A3(new_n229_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT10), .B(G99gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n220_), .B1(new_n235_), .B2(G106gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n217_), .A2(KEYINPUT65), .A3(new_n218_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n238_), .A2(KEYINPUT67), .A3(new_n212_), .A4(new_n211_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n224_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT12), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  INV_X1    g041(.A(G71gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT66), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G71gat), .ZN(new_n246_));
  INV_X1    g045(.A(G78gat), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n244_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n245_), .A2(G71gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n243_), .A2(KEYINPUT66), .ZN(new_n253_));
  OAI21_X1  g052(.A(G78gat), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n244_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT11), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n242_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(KEYINPUT11), .A3(new_n255_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n242_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n241_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n240_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G230gat), .A2(G233gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT64), .Z(new_n264_));
  OAI21_X1  g063(.A(new_n250_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n265_), .B2(new_n258_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n258_), .A2(new_n259_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G85gat), .ZN(new_n272_));
  INV_X1    g071(.A(G92gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G85gat), .A2(G92gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT9), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n212_), .A2(new_n278_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n241_), .B1(new_n268_), .B2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n268_), .A2(new_n279_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n262_), .B(new_n264_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n264_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n257_), .A2(new_n260_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n234_), .A2(new_n222_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n283_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT68), .B(G204gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G120gat), .B(G148gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(new_n293_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT69), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n295_), .A2(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(KEYINPUT69), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n300_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT97), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT95), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G197gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(G204gat), .ZN(new_n312_));
  INV_X1    g111(.A(G204gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(G197gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT21), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(KEYINPUT84), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n316_), .B(new_n317_), .C1(new_n319_), .C2(new_n312_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n310_), .A2(new_n315_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n319_), .B2(new_n312_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n308_), .A2(new_n309_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n308_), .A2(new_n309_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT21), .A4(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT23), .ZN(new_n328_));
  OR2_X1    g127(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n329_));
  NAND2_X1  g128(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n328_), .B1(new_n331_), .B2(new_n327_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n332_), .B1(G183gat), .B2(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340_));
  OR2_X1    g139(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(KEYINPUT25), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(KEYINPUT78), .ZN(new_n347_));
  OAI21_X1  g146(.A(G183gat), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n348_), .B2(KEYINPUT79), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(KEYINPUT78), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(KEYINPUT25), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n340_), .B1(new_n349_), .B2(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n354_), .A2(new_n355_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n348_), .A2(KEYINPUT79), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(KEYINPUT80), .A3(new_n359_), .A4(new_n351_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT24), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n329_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n327_), .A2(KEYINPUT23), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n335_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n357_), .A2(new_n360_), .A3(new_n363_), .A4(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n326_), .B1(new_n339_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n343_), .A2(KEYINPUT89), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n341_), .A2(new_n373_), .A3(new_n342_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n376_));
  OR3_X1    g175(.A1(new_n376_), .A2(new_n335_), .A3(new_n361_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n361_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n332_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n336_), .A2(new_n337_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n334_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n338_), .A2(KEYINPUT91), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n366_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n379_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n321_), .A2(new_n325_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n370_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT19), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n307_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n388_), .A2(new_n397_), .A3(new_n389_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n369_), .A2(new_n326_), .A3(new_n339_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n401_), .A2(KEYINPUT20), .A3(new_n395_), .A4(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n390_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n369_), .A2(new_n339_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n389_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(KEYINPUT20), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n396_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G92gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT18), .B(G64gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n388_), .A2(new_n397_), .A3(new_n389_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT20), .B(new_n402_), .C1(new_n416_), .C2(new_n398_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(new_n395_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n392_), .A2(new_n394_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(KEYINPUT27), .A3(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n401_), .A2(KEYINPUT20), .A3(new_n394_), .A4(new_n402_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n407_), .A2(new_n395_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n414_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT93), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(G155gat), .B2(G162gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT83), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(G155gat), .A3(G162gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT1), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n434_), .A2(new_n435_), .A3(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n442_), .B(KEYINPUT3), .Z(new_n446_));
  XOR2_X1   g245(.A(new_n444_), .B(KEYINPUT2), .Z(new_n447_));
  OAI211_X1 g246(.A(new_n437_), .B(new_n436_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G127gat), .B(G134gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G120gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n445_), .A2(new_n448_), .A3(new_n452_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n430_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n455_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(new_n457_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n429_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(new_n272_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT0), .B(G57gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  OR3_X1    g266(.A1(new_n460_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(KEYINPUT96), .B(new_n467_), .C1(new_n460_), .C2(new_n463_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n421_), .A2(new_n427_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n449_), .A2(KEYINPUT29), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G228gat), .A2(G233gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n389_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT29), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n326_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G78gat), .B(G106gat), .Z(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(KEYINPUT86), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n483_), .B(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(G50gat), .B1(new_n449_), .B2(KEYINPUT29), .ZN(new_n487_));
  INV_X1    g286(.A(G50gat), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n445_), .A2(new_n448_), .A3(new_n479_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT28), .B(G22gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n491_), .A3(new_n489_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n477_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT87), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n486_), .A2(new_n498_), .A3(KEYINPUT88), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n493_), .A2(new_n494_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n501_), .B1(KEYINPUT87), .B2(new_n496_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n483_), .B1(KEYINPUT86), .B2(new_n484_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n477_), .A2(new_n481_), .A3(new_n482_), .A4(new_n485_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n500_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n477_), .A2(new_n481_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(new_n484_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n508_), .A2(new_n496_), .ZN(new_n509_));
  OAI22_X1  g308(.A1(new_n499_), .A2(new_n506_), .B1(new_n509_), .B2(new_n495_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G15gat), .B(G43gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT31), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n369_), .A2(new_n513_), .A3(new_n339_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n513_), .B1(new_n369_), .B2(new_n339_), .ZN(new_n516_));
  OAI21_X1  g315(.A(G71gat), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n405_), .A2(KEYINPUT30), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(new_n243_), .A3(new_n514_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT82), .B(G99gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n512_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G227gat), .A2(G233gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n452_), .B(new_n525_), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n519_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n512_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n521_), .A3(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n526_), .B1(new_n524_), .B2(new_n531_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n510_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n526_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n522_), .A2(new_n523_), .A3(new_n512_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n530_), .B1(new_n529_), .B2(new_n521_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n495_), .B1(new_n508_), .B2(new_n496_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT88), .B1(new_n486_), .B2(new_n498_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n502_), .A2(new_n500_), .A3(new_n505_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n524_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n474_), .B1(new_n534_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n538_), .A2(new_n543_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n409_), .A2(KEYINPUT32), .A3(new_n413_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n471_), .A2(new_n549_), .A3(new_n472_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n461_), .A2(new_n430_), .A3(new_n457_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n551_), .A2(KEYINPUT94), .A3(new_n467_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n456_), .A2(new_n430_), .A3(new_n459_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT94), .B1(new_n551_), .B2(new_n467_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n420_), .A2(new_n555_), .A3(new_n424_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n469_), .B(new_n557_), .ZN(new_n558_));
  OAI22_X1  g357(.A1(new_n547_), .A2(new_n550_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n546_), .A2(new_n559_), .A3(new_n542_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n545_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G8gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT72), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT71), .B(G1gat), .ZN(new_n564_));
  INV_X1    g363(.A(G8gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G15gat), .B(G22gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n563_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G29gat), .B(G36gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n573_), .B(KEYINPUT15), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n569_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n573_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n569_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n575_), .B1(new_n574_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT77), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(KEYINPUT77), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n583_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n306_), .B1(new_n561_), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n546_), .A2(new_n559_), .A3(new_n542_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n538_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n542_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n594_), .B1(new_n597_), .B2(new_n474_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n592_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT97), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n305_), .B1(new_n593_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602_));
  XOR2_X1   g401(.A(G190gat), .B(G218gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n240_), .A2(new_n576_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT70), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(KEYINPUT35), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n279_), .A2(new_n573_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n612_), .B1(new_n610_), .B2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n602_), .B(new_n605_), .C1(new_n614_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619_));
  INV_X1    g418(.A(new_n609_), .ZN(new_n620_));
  AOI211_X1 g419(.A(new_n619_), .B(new_n620_), .C1(new_n606_), .C2(KEYINPUT70), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n606_), .B(new_n611_), .C1(new_n621_), .C2(new_n615_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n605_), .A2(new_n602_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n605_), .A2(new_n602_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .A4(new_n613_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT37), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT73), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n284_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n569_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G127gat), .B(G155gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT75), .ZN(new_n633_));
  XOR2_X1   g432(.A(G183gat), .B(G211gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT17), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n631_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n637_), .A2(KEYINPUT17), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n631_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n627_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT76), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n601_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n473_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n564_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT38), .ZN(new_n648_));
  INV_X1    g447(.A(new_n626_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n304_), .A2(new_n599_), .A3(new_n642_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(KEYINPUT98), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n598_), .B(new_n651_), .C1(KEYINPUT98), .C2(new_n650_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT99), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n473_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n654_), .ZN(G1324gat));
  NAND2_X1  g454(.A1(new_n421_), .A2(new_n427_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n652_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT39), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n645_), .A2(new_n565_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n653_), .B2(new_n546_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n546_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n645_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1326gat));
  OAI21_X1  g468(.A(G22gat), .B1(new_n653_), .B2(new_n542_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n645_), .A2(new_n672_), .A3(new_n510_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1327gat));
  NOR2_X1   g473(.A1(new_n642_), .A2(new_n626_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n601_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n646_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT37), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n626_), .B(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n598_), .A2(new_n678_), .A3(new_n679_), .A4(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n679_), .B(new_n681_), .C1(new_n545_), .C2(new_n560_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT102), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n561_), .B2(new_n627_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n642_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n304_), .A2(new_n599_), .A3(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT101), .Z(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n686_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n689_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(G29gat), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n677_), .B1(new_n693_), .B2(new_n646_), .ZN(G1328gat));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n657_), .A2(KEYINPUT103), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n657_), .A2(KEYINPUT103), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n601_), .A2(new_n695_), .A3(new_n675_), .A4(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n692_), .A2(new_n656_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G36gat), .B1(new_n702_), .B2(new_n690_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT46), .Z(G1329gat));
  NAND4_X1  g504(.A1(new_n691_), .A2(G43gat), .A3(new_n667_), .A4(new_n692_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n676_), .A2(new_n667_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G43gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n676_), .B2(new_n510_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n690_), .A2(new_n488_), .A3(new_n542_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n692_), .B2(new_n711_), .ZN(G1331gat));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n561_), .B2(new_n599_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n598_), .A2(KEYINPUT104), .A3(new_n592_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n305_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n646_), .A3(new_n644_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n598_), .A2(new_n592_), .A3(new_n626_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n305_), .A2(new_n642_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n473_), .A2(new_n718_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n717_), .A2(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1332gat));
  INV_X1    g522(.A(G64gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n721_), .B2(new_n699_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT48), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n716_), .A2(new_n644_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n699_), .A2(new_n724_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(G1333gat));
  AOI21_X1  g528(.A(new_n243_), .B1(new_n721_), .B2(new_n667_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT49), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n667_), .A2(new_n243_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n727_), .B2(new_n732_), .ZN(G1334gat));
  AOI21_X1  g532(.A(new_n247_), .B1(new_n721_), .B2(new_n510_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n542_), .A2(G78gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT106), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n727_), .B2(new_n738_), .ZN(G1335gat));
  NOR3_X1   g538(.A1(new_n304_), .A2(new_n599_), .A3(new_n642_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n686_), .A2(new_n740_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n741_), .A2(new_n272_), .A3(new_n473_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n716_), .A2(KEYINPUT107), .A3(new_n675_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n714_), .A2(new_n715_), .A3(new_n305_), .A4(new_n675_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n646_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT108), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT108), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n742_), .B1(new_n749_), .B2(new_n750_), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n741_), .A2(new_n273_), .A3(new_n698_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n747_), .A2(new_n656_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n273_), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n217_), .A3(new_n667_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G99gat), .B1(new_n741_), .B2(new_n546_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n747_), .A2(KEYINPUT109), .A3(new_n217_), .A4(new_n667_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT51), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n757_), .A2(new_n759_), .A3(new_n762_), .A4(new_n758_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1338gat));
  XNOR2_X1  g563(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n686_), .A2(new_n510_), .A3(new_n740_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(G106gat), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT110), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n775_), .ZN(new_n776_));
  AOI211_X1 g575(.A(G106gat), .B(new_n542_), .C1(new_n743_), .C2(new_n746_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n765_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n765_), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n777_), .C1(new_n770_), .C2(new_n775_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  INV_X1    g581(.A(new_n300_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n295_), .A2(new_n296_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n592_), .B(new_n642_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n304_), .A2(KEYINPUT112), .A3(new_n592_), .A4(new_n642_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n627_), .A3(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT114), .Z(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n583_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n574_), .A2(new_n581_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n575_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n574_), .A2(new_n577_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n801_), .B(new_n588_), .C1(new_n575_), .C2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n301_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n282_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n262_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n283_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT12), .B1(new_n284_), .B2(new_n285_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n284_), .A2(new_n285_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(KEYINPUT55), .A3(new_n264_), .A4(new_n262_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(new_n809_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT115), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n807_), .A2(new_n813_), .A3(new_n809_), .A4(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n293_), .A4(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n293_), .A3(new_n817_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n820_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n818_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n592_), .A2(new_n294_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n805_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n798_), .B1(new_n826_), .B2(new_n649_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n825_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n819_), .A2(new_n821_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT116), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n818_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT57), .B(new_n626_), .C1(new_n833_), .C2(new_n805_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n799_), .A2(new_n295_), .A3(new_n803_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n829_), .B2(new_n818_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n649_), .A2(KEYINPUT37), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n626_), .A2(new_n680_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(KEYINPUT58), .A2(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n829_), .A2(new_n818_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n836_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n835_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n841_), .A2(KEYINPUT58), .A3(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n681_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n844_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n837_), .A2(new_n849_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n848_), .A2(KEYINPUT118), .A3(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n827_), .B(new_n834_), .C1(new_n846_), .C2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n797_), .B1(new_n852_), .B2(new_n687_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n544_), .A2(new_n473_), .A3(new_n656_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n599_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n840_), .A2(new_n845_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n827_), .A2(new_n834_), .A3(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n860_), .A2(new_n687_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n797_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n854_), .A2(new_n858_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n856_), .A2(new_n858_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n599_), .A2(G113gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n857_), .B1(new_n865_), .B2(new_n866_), .ZN(G1340gat));
  OR3_X1    g666(.A1(new_n864_), .A2(KEYINPUT119), .A3(new_n304_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n864_), .B2(new_n304_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(G120gat), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n856_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n856_), .B2(new_n642_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n642_), .A2(G127gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n865_), .B2(new_n876_), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n856_), .B2(new_n649_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n681_), .A2(G134gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n865_), .B2(new_n879_), .ZN(G1343gat));
  NOR4_X1   g679(.A1(new_n853_), .A2(new_n473_), .A3(new_n534_), .A4(new_n699_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n599_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT120), .B(G141gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n305_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n642_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  AOI21_X1  g688(.A(G162gat), .B1(new_n881_), .B2(new_n649_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n681_), .A2(G162gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n881_), .B2(new_n891_), .ZN(G1347gat));
  NOR3_X1   g691(.A1(new_n698_), .A2(new_n646_), .A3(new_n546_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n542_), .B(new_n893_), .C1(new_n861_), .C2(new_n797_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G169gat), .B1(new_n894_), .B2(new_n592_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(KEYINPUT121), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(KEYINPUT121), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(KEYINPUT62), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(KEYINPUT121), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n894_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n599_), .A3(new_n336_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(new_n900_), .A3(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n901_), .B2(new_n305_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n893_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n826_), .A2(new_n649_), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n848_), .B2(new_n850_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n840_), .A2(new_n835_), .A3(new_n845_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(KEYINPUT57), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n642_), .B1(new_n909_), .B2(new_n827_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT122), .B(new_n542_), .C1(new_n910_), .C2(new_n797_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n853_), .B2(new_n510_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n905_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n304_), .A2(new_n337_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n904_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NOR3_X1   g715(.A1(new_n894_), .A2(new_n687_), .A3(new_n372_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n913_), .ZN(new_n919_));
  AND4_X1   g718(.A1(new_n918_), .A2(new_n919_), .A3(new_n642_), .A4(new_n893_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n914_), .B2(new_n642_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n917_), .B1(new_n922_), .B2(new_n350_), .ZN(G1350gat));
  NAND4_X1  g722(.A1(new_n901_), .A2(new_n649_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G190gat), .B1(new_n894_), .B2(new_n627_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT124), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n596_), .A2(new_n473_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n853_), .B1(KEYINPUT125), .B2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n928_), .A2(KEYINPUT125), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n698_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n592_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n311_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n304_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n313_), .ZN(G1353gat));
  XNOR2_X1  g735(.A(KEYINPUT63), .B(G211gat), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n929_), .A2(new_n642_), .A3(new_n931_), .A4(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n932_), .A2(new_n687_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n938_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT126), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n943_), .B(new_n938_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n944_), .ZN(G1354gat));
  OAI21_X1  g744(.A(G218gat), .B1(new_n932_), .B2(new_n627_), .ZN(new_n946_));
  INV_X1    g745(.A(G218gat), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n929_), .A2(new_n947_), .A3(new_n649_), .A4(new_n931_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(KEYINPUT127), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n946_), .A2(new_n951_), .A3(new_n948_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(G1355gat));
endmodule


