//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n970_, new_n971_,
    new_n972_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n988_, new_n990_, new_n991_, new_n992_, new_n994_,
    new_n995_, new_n996_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(G197gat), .B(G204gat), .Z(new_n209_));
  OAI211_X1 g008(.A(KEYINPUT21), .B(new_n208_), .C1(new_n209_), .C2(KEYINPUT87), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n205_), .A2(new_n204_), .ZN(new_n211_));
  AOI22_X1  g010(.A1(new_n206_), .A2(new_n210_), .B1(new_n203_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G190gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT77), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G183gat), .A3(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT23), .ZN(new_n233_));
  NOR3_X1   g032(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT92), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(new_n232_), .B2(KEYINPUT23), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT92), .A3(new_n235_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n227_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n225_), .ZN(new_n244_));
  INV_X1    g043(.A(G169gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT22), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G169gat), .ZN(new_n248_));
  INV_X1    g047(.A(G176gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n228_), .A2(KEYINPUT76), .A3(KEYINPUT23), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT76), .B1(new_n228_), .B2(KEYINPUT23), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT23), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n232_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n214_), .A2(new_n218_), .ZN(new_n258_));
  AOI211_X1 g057(.A(new_n244_), .B(new_n251_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n213_), .B1(new_n243_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT93), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n227_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n222_), .A2(new_n226_), .A3(KEYINPUT75), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n235_), .A3(new_n257_), .A4(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n244_), .B1(new_n250_), .B2(KEYINPUT78), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n246_), .A2(new_n248_), .A3(new_n268_), .A4(new_n249_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n250_), .A2(KEYINPUT78), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(new_n266_), .A3(new_n225_), .A4(new_n269_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n233_), .A2(new_n258_), .A3(new_n237_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n265_), .B(new_n212_), .C1(new_n270_), .C2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n275_), .A2(KEYINPUT20), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT91), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT25), .B(G183gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G190gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n281_), .A2(new_n282_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT92), .B1(new_n241_), .B2(new_n235_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n255_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n285_));
  NOR4_X1   g084(.A1(new_n285_), .A2(new_n239_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n283_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n257_), .A2(new_n258_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n251_), .A2(new_n244_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT93), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n213_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n261_), .A2(new_n276_), .A3(new_n280_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n257_), .A2(new_n264_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n235_), .B1(new_n283_), .B2(KEYINPUT75), .ZN(new_n296_));
  OAI22_X1  g095(.A1(new_n274_), .A2(new_n270_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n213_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n290_), .A3(new_n212_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(KEYINPUT20), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n280_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G8gat), .B(G36gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n294_), .A2(new_n302_), .A3(new_n309_), .ZN(new_n310_));
  AND4_X1   g109(.A1(KEYINPUT20), .A2(new_n298_), .A3(new_n280_), .A4(new_n299_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n261_), .A2(new_n276_), .A3(new_n293_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n301_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n313_), .B2(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(G155gat), .ZN(new_n316_));
  INV_X1    g115(.A(G162gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(KEYINPUT84), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n319_), .B1(G155gat), .B2(G162gat), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n318_), .A2(new_n320_), .B1(G155gat), .B2(G162gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n323_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n321_), .B1(new_n327_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n322_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(new_n328_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n318_), .A2(new_n320_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT1), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G134gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G127gat), .ZN(new_n345_));
  INV_X1    g144(.A(G127gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G134gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n343_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n346_), .A2(G134gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n344_), .A2(G127gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT81), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(new_n342_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n334_), .A2(new_n341_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n315_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n337_), .A2(new_n339_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(new_n323_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n336_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n339_), .B(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n337_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n360_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n334_), .A2(new_n341_), .A3(new_n356_), .A4(new_n351_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT4), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n359_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT96), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  NAND3_X1  g177(.A1(new_n370_), .A2(new_n371_), .A3(new_n315_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT96), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n359_), .A2(new_n372_), .A3(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n374_), .A2(new_n378_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT97), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n381_), .A2(new_n379_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n385_), .A2(KEYINPUT97), .A3(new_n378_), .A4(new_n374_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n378_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n379_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n380_), .B1(new_n359_), .B2(new_n372_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n314_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n292_), .B1(new_n291_), .B2(new_n213_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n275_), .A2(KEYINPUT20), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n280_), .B1(new_n395_), .B2(new_n293_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n307_), .B1(new_n396_), .B2(new_n311_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n312_), .A2(new_n301_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n311_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n308_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(KEYINPUT95), .B(new_n307_), .C1(new_n396_), .C2(new_n311_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n382_), .A2(KEYINPUT33), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n385_), .A2(new_n406_), .A3(new_n378_), .A4(new_n374_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n334_), .A2(new_n341_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n372_), .A2(new_n315_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n370_), .A2(new_n371_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n411_), .B(new_n387_), .C1(new_n412_), .C2(new_n315_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n392_), .B1(new_n404_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT86), .B1(new_n419_), .B2(new_n212_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n213_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n420_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n409_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G22gat), .B(G50gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n427_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n438_), .B(KEYINPUT88), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n425_), .A2(new_n426_), .A3(new_n443_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT89), .B1(new_n434_), .B2(new_n436_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n427_), .A2(new_n446_), .A3(new_n442_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n441_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n202_), .B1(new_n416_), .B2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n414_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT98), .B(new_n449_), .C1(new_n452_), .C2(new_n392_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n449_), .A2(new_n391_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT27), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n402_), .A2(new_n403_), .A3(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n294_), .A2(new_n302_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n401_), .B(KEYINPUT27), .C1(new_n308_), .C2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n454_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(new_n453_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(G71gat), .Z(new_n462_));
  INV_X1    g261(.A(G99gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n297_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT83), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n297_), .A2(new_n464_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT80), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT30), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(new_n360_), .ZN(new_n474_));
  OR3_X1    g273(.A1(new_n469_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n474_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n391_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n456_), .A2(new_n449_), .A3(new_n458_), .A4(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT99), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n460_), .A2(new_n478_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT100), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G169gat), .B(G197gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G8gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT72), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(KEYINPUT72), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493_));
  INV_X1    g292(.A(G1gat), .ZN(new_n494_));
  INV_X1    g293(.A(G8gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n490_), .A2(new_n496_), .A3(new_n493_), .A4(new_n491_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n499_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n503_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(G229gat), .B(G233gat), .C1(new_n504_), .C2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n503_), .B(KEYINPUT15), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n503_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT73), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n488_), .B1(new_n515_), .B2(KEYINPUT74), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n517_));
  INV_X1    g316(.A(new_n488_), .ZN(new_n518_));
  AOI211_X1 g317(.A(new_n517_), .B(new_n518_), .C1(new_n508_), .C2(new_n514_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR3_X1   g320(.A1(new_n484_), .A2(new_n485_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n485_), .B1(new_n484_), .B2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G85gat), .B(G92gat), .Z(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(KEYINPUT9), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT10), .B(G99gat), .Z(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT64), .B(G85gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(G92gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n463_), .A3(new_n532_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n529_), .B1(new_n528_), .B2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(KEYINPUT8), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(KEYINPUT8), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT66), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT66), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n547_), .B(new_n537_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n509_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT70), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n546_), .A2(new_n551_), .A3(new_n509_), .A4(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT34), .ZN(new_n555_));
  OAI22_X1  g354(.A1(new_n545_), .A2(new_n506_), .B1(KEYINPUT35), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n555_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT35), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT71), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n553_), .A2(new_n564_), .A3(new_n557_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n553_), .B2(new_n557_), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n561_), .B(new_n556_), .C1(new_n550_), .C2(new_n552_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT71), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n572_), .B(KEYINPUT36), .Z(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n562_), .A2(new_n575_), .A3(new_n565_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT37), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n573_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n578_), .A3(KEYINPUT37), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n505_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G71gat), .B(G78gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT11), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(KEYINPUT11), .ZN(new_n587_));
  INV_X1    g386(.A(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n584_), .A2(KEYINPUT11), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n586_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n583_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT17), .ZN(new_n599_));
  AND2_X1   g398(.A1(KEYINPUT67), .A2(KEYINPUT17), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n593_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n581_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n537_), .B(new_n591_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n545_), .A2(new_n592_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT12), .B1(new_n591_), .B2(KEYINPUT67), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(KEYINPUT67), .B2(new_n591_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n611_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n612_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT65), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n610_), .B1(new_n618_), .B2(new_n607_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n608_), .A2(KEYINPUT65), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT5), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n616_), .A2(new_n621_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(KEYINPUT68), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT68), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n631_), .A3(new_n626_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n630_), .A2(KEYINPUT13), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT13), .B1(new_n630_), .B2(new_n632_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT69), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT69), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n606_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n525_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n525_), .A2(KEYINPUT101), .A3(new_n640_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n643_), .A2(new_n494_), .A3(new_n391_), .A4(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT102), .B1(new_n639_), .B2(new_n521_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n636_), .A2(new_n649_), .A3(new_n520_), .A4(new_n638_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n605_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n460_), .A2(new_n478_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n483_), .A2(new_n482_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n574_), .A2(new_n576_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT103), .B1(new_n484_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n651_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n391_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G1gat), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n645_), .A2(new_n646_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n647_), .A2(new_n663_), .A3(new_n664_), .ZN(G1324gat));
  AND2_X1   g464(.A1(new_n456_), .A2(new_n458_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(G8gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n643_), .A2(new_n644_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  INV_X1    g468(.A(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n660_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n671_), .B2(G8gat), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT39), .B(new_n495_), .C1(new_n660_), .C2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n668_), .B(KEYINPUT40), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1325gat));
  NAND2_X1  g477(.A1(new_n643_), .A2(new_n644_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n478_), .A2(G15gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n660_), .A2(new_n477_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n679_), .A2(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1326gat));
  INV_X1    g483(.A(G22gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n450_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n660_), .A2(new_n450_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(G22gat), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT42), .B(new_n685_), .C1(new_n660_), .C2(new_n450_), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n679_), .A2(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(G1327gat));
  NOR2_X1   g490(.A1(new_n656_), .A2(new_n605_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n639_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n525_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G29gat), .B1(new_n696_), .B2(new_n391_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT37), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n656_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n579_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n484_), .B2(new_n581_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n581_), .B2(KEYINPUT104), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n449_), .B1(new_n452_), .B2(new_n392_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n202_), .A2(new_n706_), .B1(new_n666_), .B2(new_n454_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n477_), .B1(new_n707_), .B2(new_n453_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n483_), .A2(new_n482_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n705_), .B(new_n701_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n704_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n605_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n648_), .A2(new_n712_), .A3(new_n650_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT44), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n716_), .B(new_n713_), .C1(new_n704_), .C2(new_n710_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n391_), .A2(G29gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n697_), .B1(new_n718_), .B2(new_n719_), .ZN(G1328gat));
  INV_X1    g519(.A(new_n715_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n711_), .A2(KEYINPUT44), .A3(new_n714_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n670_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n666_), .A2(G36gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT100), .B1(new_n654_), .B2(new_n520_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n694_), .B(new_n726_), .C1(new_n727_), .C2(new_n522_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT106), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n728_), .A2(new_n731_), .B1(KEYINPUT107), .B2(KEYINPUT46), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n728_), .A2(new_n731_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n724_), .A2(new_n725_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n725_), .B1(new_n724_), .B2(new_n734_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n695_), .B2(new_n478_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n478_), .A2(new_n738_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n715_), .A2(new_n717_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NOR4_X1   g543(.A1(new_n715_), .A2(new_n717_), .A3(KEYINPUT108), .A4(new_n741_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT47), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n718_), .A2(new_n740_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT108), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n742_), .A2(new_n743_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .A4(new_n739_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n746_), .A2(new_n751_), .ZN(G1330gat));
  NOR3_X1   g551(.A1(new_n715_), .A2(new_n717_), .A3(new_n449_), .ZN(new_n753_));
  INV_X1    g552(.A(G50gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n450_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT109), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n753_), .A2(new_n754_), .B1(new_n695_), .B2(new_n756_), .ZN(G1331gat));
  NAND2_X1  g556(.A1(new_n657_), .A2(new_n659_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n639_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n521_), .A2(new_n605_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G57gat), .B1(new_n762_), .B2(new_n662_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n484_), .A2(new_n520_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n759_), .A2(new_n606_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n766_), .A2(G57gat), .A3(new_n662_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n767_), .ZN(G1332gat));
  INV_X1    g567(.A(new_n766_), .ZN(new_n769_));
  INV_X1    g568(.A(G64gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n670_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772_));
  INV_X1    g571(.A(new_n762_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n670_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n774_), .B2(G64gat), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT48), .B(new_n770_), .C1(new_n773_), .C2(new_n670_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n775_), .B2(new_n776_), .ZN(G1333gat));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n477_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G71gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G71gat), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n478_), .A2(G71gat), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT110), .ZN(new_n783_));
  OAI22_X1  g582(.A1(new_n780_), .A2(new_n781_), .B1(new_n766_), .B2(new_n783_), .ZN(G1334gat));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n769_), .A2(new_n785_), .A3(new_n450_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n773_), .A2(new_n450_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G78gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT50), .B(new_n785_), .C1(new_n773_), .C2(new_n450_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1335gat));
  NAND3_X1  g590(.A1(new_n764_), .A2(new_n639_), .A3(new_n692_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(new_n662_), .ZN(new_n793_));
  INV_X1    g592(.A(G85gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n639_), .A2(new_n521_), .A3(new_n712_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n704_), .B2(new_n710_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n391_), .A2(new_n534_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT111), .Z(new_n798_));
  AOI22_X1  g597(.A1(new_n793_), .A2(new_n794_), .B1(new_n796_), .B2(new_n798_), .ZN(G1336gat));
  AND2_X1   g598(.A1(new_n796_), .A2(new_n670_), .ZN(new_n800_));
  INV_X1    g599(.A(G92gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n670_), .A2(new_n801_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n800_), .A2(new_n801_), .B1(new_n792_), .B2(new_n802_), .ZN(G1337gat));
  AND2_X1   g602(.A1(new_n796_), .A2(new_n477_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n477_), .A2(new_n531_), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n804_), .A2(new_n463_), .B1(new_n792_), .B2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT113), .B(new_n532_), .C1(new_n796_), .C2(new_n450_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810_));
  INV_X1    g609(.A(new_n795_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n705_), .B1(new_n654_), .B2(new_n701_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n484_), .A2(new_n581_), .A3(new_n703_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n450_), .B(new_n811_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n814_), .B2(G106gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n808_), .B1(new_n809_), .B2(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n449_), .B(new_n795_), .C1(new_n704_), .C2(new_n710_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n817_), .B2(new_n532_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n810_), .A3(G106gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT52), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n450_), .A2(new_n532_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n792_), .A2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT112), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT53), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n816_), .A2(new_n820_), .A3(new_n826_), .A4(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1339gat));
  NOR2_X1   g627(.A1(new_n635_), .A2(new_n760_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n829_), .A2(new_n581_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n829_), .B2(new_n581_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n612_), .B1(new_n611_), .B2(new_n615_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n616_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n611_), .A2(new_n615_), .A3(KEYINPUT55), .A4(new_n612_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n626_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n520_), .A2(new_n629_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n838_), .B2(new_n626_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n843_), .B(new_n628_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n841_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n513_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n513_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n510_), .A2(new_n511_), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  MUX2_X1   g650(.A(new_n851_), .B(new_n515_), .S(new_n488_), .Z(new_n852_));
  NAND3_X1  g651(.A1(new_n630_), .A2(new_n632_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n630_), .A2(KEYINPUT115), .A3(new_n632_), .A4(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n656_), .B1(new_n847_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n861_));
  NAND2_X1  g660(.A1(new_n852_), .A2(new_n629_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n845_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n862_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n864_), .B(KEYINPUT58), .C1(new_n842_), .C2(new_n844_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT117), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n838_), .A2(new_n626_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n843_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n838_), .A2(KEYINPUT56), .A3(new_n626_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(KEYINPUT58), .A4(new_n864_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n701_), .A2(new_n863_), .A3(new_n866_), .A4(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n842_), .A2(new_n844_), .A3(KEYINPUT114), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n855_), .B(new_n856_), .C1(new_n874_), .C2(new_n841_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT57), .A3(new_n656_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n860_), .A2(new_n873_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n833_), .B1(new_n877_), .B2(new_n712_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n670_), .A2(new_n450_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n478_), .A2(new_n662_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n872_), .A2(new_n866_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n862_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n861_), .ZN(new_n887_));
  OAI22_X1  g686(.A1(new_n577_), .A2(new_n580_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n885_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n875_), .B2(new_n656_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n884_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n860_), .A2(new_n873_), .A3(KEYINPUT118), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n876_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n833_), .B1(new_n893_), .B2(new_n712_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n881_), .A2(KEYINPUT59), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  OAI22_X1  g695(.A1(new_n882_), .A2(new_n883_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G113gat), .B1(new_n897_), .B2(new_n521_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n882_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n521_), .A2(G113gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1340gat));
  OAI21_X1  g700(.A(G120gat), .B1(new_n897_), .B2(new_n759_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903_));
  AOI21_X1  g702(.A(G120gat), .B1(new_n639_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT119), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(new_n903_), .B2(G120gat), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n882_), .B(new_n905_), .C1(new_n904_), .C2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n902_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT120), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n902_), .A2(new_n911_), .A3(new_n908_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1341gat));
  OAI21_X1  g712(.A(G127gat), .B1(new_n897_), .B2(new_n712_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n882_), .A2(new_n346_), .A3(new_n605_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1342gat));
  AOI21_X1  g715(.A(G134gat), .B1(new_n882_), .B2(new_n658_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n897_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT121), .B(G134gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n581_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n918_), .B2(new_n920_), .ZN(G1343gat));
  NAND2_X1  g720(.A1(new_n877_), .A2(new_n712_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n833_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n450_), .A2(new_n478_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n670_), .A2(new_n662_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n521_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT122), .B(G141gat), .Z(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1344gat));
  INV_X1    g729(.A(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n639_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g732(.A1(new_n927_), .A2(new_n712_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n927_), .B2(new_n581_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n658_), .A2(new_n317_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n927_), .B2(new_n940_), .ZN(G1347gat));
  NAND2_X1  g740(.A1(new_n670_), .A2(new_n479_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n450_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n893_), .A2(new_n712_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n923_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n245_), .B1(new_n946_), .B2(new_n520_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n948_));
  OAI21_X1  g747(.A(KEYINPUT125), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n894_), .A2(new_n521_), .A3(new_n944_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n950_), .B(KEYINPUT62), .C1(new_n951_), .C2(new_n245_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n876_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n860_), .A2(new_n873_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n884_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n605_), .B1(new_n955_), .B2(new_n892_), .ZN(new_n956_));
  OAI211_X1 g755(.A(new_n520_), .B(new_n943_), .C1(new_n956_), .C2(new_n833_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n957_), .A2(new_n948_), .A3(G169gat), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n957_), .A2(KEYINPUT124), .A3(new_n948_), .A4(G169gat), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n949_), .A2(new_n952_), .A3(new_n960_), .A4(new_n961_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n951_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1348gat));
  AOI21_X1  g763(.A(G176gat), .B1(new_n946_), .B2(new_n639_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n924_), .A2(new_n449_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n759_), .A2(new_n249_), .A3(new_n942_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n965_), .B1(new_n967_), .B2(new_n968_), .ZN(G1349gat));
  INV_X1    g768(.A(new_n946_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n970_), .A2(new_n281_), .A3(new_n712_), .ZN(new_n971_));
  OR3_X1    g770(.A1(new_n966_), .A2(new_n712_), .A3(new_n942_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(new_n214_), .B2(new_n972_), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n946_), .A2(new_n282_), .A3(new_n658_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n970_), .A2(new_n581_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n218_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(KEYINPUT126), .ZN(new_n977_));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978_));
  OAI211_X1 g777(.A(new_n978_), .B(new_n974_), .C1(new_n975_), .C2(new_n218_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n977_), .A2(new_n979_), .ZN(G1351gat));
  NOR3_X1   g779(.A1(new_n925_), .A2(new_n666_), .A3(new_n391_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n924_), .A2(new_n981_), .ZN(new_n982_));
  OR2_X1    g781(.A1(new_n982_), .A2(KEYINPUT127), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n982_), .A2(KEYINPUT127), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n985_), .A2(new_n520_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n986_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g786(.A1(new_n985_), .A2(new_n639_), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n988_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g788(.A(KEYINPUT63), .B(G211gat), .C1(new_n985_), .C2(new_n605_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(KEYINPUT63), .B(G211gat), .ZN(new_n991_));
  AOI211_X1 g790(.A(new_n712_), .B(new_n991_), .C1(new_n983_), .C2(new_n984_), .ZN(new_n992_));
  NOR2_X1   g791(.A1(new_n990_), .A2(new_n992_), .ZN(G1354gat));
  INV_X1    g792(.A(G218gat), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n985_), .A2(new_n994_), .A3(new_n658_), .ZN(new_n995_));
  AOI21_X1  g794(.A(new_n581_), .B1(new_n983_), .B2(new_n984_), .ZN(new_n996_));
  OAI21_X1  g795(.A(new_n995_), .B1(new_n994_), .B2(new_n996_), .ZN(G1355gat));
endmodule


