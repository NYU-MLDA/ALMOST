//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(KEYINPUT88), .B2(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(KEYINPUT88), .B2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  AOI21_X1  g006(.A(G176gat), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n205_), .B(new_n208_), .C1(new_n207_), .C2(new_n206_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT89), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT83), .B(G183gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT23), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n212_), .B1(new_n214_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n210_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n219_), .B(KEYINPUT86), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n223_), .A2(new_n217_), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n202_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(KEYINPUT24), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n213_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n216_), .B2(KEYINPUT26), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(G183gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n233_), .A2(new_n235_), .A3(new_n236_), .A4(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n229_), .B1(new_n231_), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT85), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT85), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n228_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n222_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G99gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT90), .B(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  XOR2_X1   g046(.A(G127gat), .B(G134gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT91), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT31), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n247_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(G15gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT30), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT92), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n260_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT97), .B(G197gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(KEYINPUT21), .A3(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n266_), .A2(G204gat), .ZN(new_n271_));
  INV_X1    g070(.A(G197gat), .ZN(new_n272_));
  INV_X1    g071(.A(G204gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT21), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n268_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n270_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n227_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n215_), .A2(KEYINPUT25), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n236_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n234_), .A2(G190gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n237_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n278_), .A2(new_n229_), .A3(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n203_), .A2(G169gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n206_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n212_), .B1(new_n286_), .B2(new_n225_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(KEYINPUT98), .B(new_n287_), .C1(new_n224_), .C2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n224_), .B2(new_n288_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT98), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n284_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n277_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n222_), .B2(new_n242_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT19), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT20), .ZN(new_n299_));
  OR3_X1    g098(.A1(new_n293_), .A2(new_n295_), .A3(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n222_), .A2(new_n294_), .A3(new_n242_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n283_), .B1(new_n292_), .B2(new_n289_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n301_), .B(KEYINPUT20), .C1(new_n302_), .C2(new_n294_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n297_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G8gat), .B(G36gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT100), .ZN(new_n306_));
  XOR2_X1   g105(.A(G64gat), .B(G92gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  AND3_X1   g109(.A1(new_n300_), .A2(new_n304_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n310_), .B(KEYINPUT104), .ZN(new_n314_));
  INV_X1    g113(.A(new_n290_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT20), .B1(new_n284_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n297_), .B1(new_n295_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n317_), .B1(new_n303_), .B2(new_n297_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n310_), .B1(new_n300_), .B2(new_n304_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n311_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n329_));
  OR2_X1    g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT1), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n335_), .A2(KEYINPUT3), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(KEYINPUT3), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n331_), .A2(new_n332_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT96), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(KEYINPUT96), .A3(new_n344_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n254_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT101), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n337_), .A2(new_n344_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT102), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n349_), .A2(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT4), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n349_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n352_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n328_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n355_), .B(KEYINPUT102), .ZN(new_n364_));
  INV_X1    g163(.A(new_n361_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n351_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n327_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n277_), .B1(new_n353_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G228gat), .A3(G233gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n347_), .A2(new_n348_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n277_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n372_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G78gat), .B(G106gat), .Z(new_n378_));
  OR2_X1    g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT28), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n373_), .B2(new_n370_), .ZN(new_n381_));
  AOI211_X1 g180(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n347_), .C2(new_n348_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G22gat), .B(G50gat), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n378_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n379_), .A2(new_n385_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n377_), .A2(new_n378_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n377_), .A2(new_n378_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n386_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n389_), .A2(new_n390_), .B1(new_n391_), .B2(new_n384_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  NOR4_X1   g192(.A1(new_n264_), .A2(new_n323_), .A3(new_n369_), .A4(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n310_), .A2(KEYINPUT32), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n300_), .A2(new_n304_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n318_), .A2(KEYINPUT32), .A3(new_n310_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT103), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n397_), .A2(KEYINPUT103), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n369_), .A2(new_n396_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n368_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n311_), .A2(new_n321_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n352_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(new_n328_), .C1(new_n352_), .C2(new_n358_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n364_), .A2(KEYINPUT33), .A3(new_n327_), .A4(new_n367_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n393_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n323_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n363_), .A2(new_n368_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n393_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n261_), .A2(KEYINPUT93), .A3(new_n262_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT93), .B1(new_n261_), .B2(new_n262_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n394_), .B1(new_n414_), .B2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G113gat), .B(G141gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT81), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT82), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G169gat), .B(G197gat), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G8gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G15gat), .B(G22gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT76), .B(G1gat), .ZN(new_n429_));
  INV_X1    g228(.A(G8gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT77), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n435_), .B(new_n428_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n427_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G29gat), .B(G36gat), .Z(new_n439_));
  XOR2_X1   g238(.A(G43gat), .B(G50gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT15), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n434_), .A2(new_n436_), .A3(new_n427_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n441_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n443_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(new_n437_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G229gat), .A2(G233gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n441_), .B(KEYINPUT79), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n438_), .A2(new_n452_), .A3(new_n443_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n449_), .B1(new_n453_), .B2(new_n448_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT80), .B(new_n426_), .C1(new_n451_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n454_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n426_), .A2(KEYINPUT80), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(new_n450_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n419_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G190gat), .B(G218gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G134gat), .B(G162gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT36), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OR3_X1    g269(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT66), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n474_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .A4(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT67), .ZN(new_n478_));
  OR2_X1    g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n477_), .A2(KEYINPUT67), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n476_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n478_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n485_));
  INV_X1    g284(.A(G85gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n487_));
  AND2_X1   g286(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n479_), .A2(KEYINPUT9), .A3(new_n480_), .ZN(new_n491_));
  OR2_X1    g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .A4(new_n470_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n484_), .A2(new_n485_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n441_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT75), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G232gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n500_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n468_), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n471_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n473_), .A2(new_n475_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n483_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n478_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n476_), .A2(new_n478_), .A3(new_n483_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(KEYINPUT70), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n496_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT73), .B1(new_n520_), .B2(new_n442_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n497_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT73), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n441_), .B(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n522_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n507_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n503_), .A2(new_n504_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n520_), .A2(KEYINPUT73), .A3(new_n442_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n523_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n528_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n507_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n465_), .B1(new_n529_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n464_), .A2(KEYINPUT36), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n533_), .B1(new_n532_), .B2(new_n507_), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n528_), .B(new_n506_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n537_), .B1(new_n540_), .B2(KEYINPUT74), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n529_), .A2(KEYINPUT74), .A3(new_n534_), .A4(new_n537_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n536_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT37), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n529_), .A2(KEYINPUT74), .A3(new_n534_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n535_), .B1(new_n548_), .B2(new_n542_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(G64gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(G57gat), .ZN(new_n553_));
  INV_X1    g352(.A(G57gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G64gat), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n553_), .A2(new_n555_), .A3(KEYINPUT68), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT68), .B1(new_n553_), .B2(new_n555_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT11), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n554_), .A2(G64gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n552_), .A2(G57gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT11), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n553_), .A2(new_n555_), .A3(KEYINPUT68), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT11), .B(new_n566_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n438_), .A2(new_n443_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(KEYINPUT71), .A2(KEYINPUT78), .ZN(new_n580_));
  AND2_X1   g379(.A1(KEYINPUT71), .A2(KEYINPUT78), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n579_), .B(KEYINPUT17), .C1(new_n580_), .C2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n582_), .B1(KEYINPUT17), .B2(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n574_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n570_), .A2(KEYINPUT71), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT71), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n568_), .A2(new_n588_), .A3(new_n569_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n587_), .A2(KEYINPUT12), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n570_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n516_), .A2(new_n496_), .A3(new_n517_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT12), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n590_), .A2(new_n520_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT64), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n498_), .A2(new_n570_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n594_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT69), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT5), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  NAND2_X1  g407(.A1(new_n604_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n598_), .A2(new_n602_), .A3(new_n603_), .A4(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n609_), .A2(KEYINPUT13), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT13), .B1(new_n609_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n545_), .A2(new_n551_), .A3(new_n586_), .A4(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n461_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT105), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n461_), .A2(KEYINPUT105), .A3(new_n616_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n369_), .A2(new_n429_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT38), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n549_), .B(KEYINPUT106), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n419_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n614_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n586_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n626_), .A2(new_n460_), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n412_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT38), .B1(new_n621_), .B2(new_n622_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT107), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT107), .B(KEYINPUT38), .C1(new_n621_), .C2(new_n622_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n634_), .B2(new_n635_), .ZN(G1324gat));
  XNOR2_X1  g435(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n625_), .A2(new_n323_), .A3(new_n628_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n638_), .B2(G8gat), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n619_), .A2(new_n430_), .A3(new_n323_), .A4(new_n620_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n637_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n644_), .B(new_n637_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1325gat));
  NAND3_X1  g447(.A1(new_n625_), .A2(new_n417_), .A3(new_n628_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G15gat), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT109), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT109), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(KEYINPUT41), .A3(new_n652_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n617_), .A2(G15gat), .A3(new_n418_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n629_), .B2(new_n409_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n409_), .A2(G22gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n617_), .B2(new_n661_), .ZN(G1327gat));
  NOR3_X1   g461(.A1(new_n626_), .A2(new_n549_), .A3(new_n586_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n461_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G29gat), .B1(new_n665_), .B2(new_n369_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n549_), .A2(new_n550_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT37), .B(new_n535_), .C1(new_n548_), .C2(new_n542_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(KEYINPUT111), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n417_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n670_), .B(new_n673_), .C1(new_n674_), .C2(new_n394_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n393_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n412_), .A2(new_n393_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n323_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n418_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n394_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n669_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n675_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n614_), .A2(new_n459_), .A3(new_n627_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT110), .Z(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT44), .B1(new_n683_), .B2(new_n686_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n369_), .A2(G29gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n666_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n411_), .A2(KEYINPUT112), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n320_), .A2(KEYINPUT112), .A3(new_n322_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n461_), .A2(new_n692_), .A3(new_n663_), .A4(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n687_), .A2(new_n688_), .A3(new_n411_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n692_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI221_X1 g501(.A(new_n698_), .B1(KEYINPUT113), .B2(KEYINPUT46), .C1(new_n699_), .C2(new_n692_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n264_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n689_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n664_), .B2(new_n418_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n665_), .B2(new_n393_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n393_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n689_), .B2(new_n714_), .ZN(G1331gat));
  NAND4_X1  g514(.A1(new_n625_), .A2(new_n460_), .A3(new_n586_), .A4(new_n626_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n412_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n419_), .A2(new_n459_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n667_), .A2(new_n668_), .A3(new_n627_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n626_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n369_), .A2(new_n554_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n716_), .B2(new_n695_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n695_), .A2(G64gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT115), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n720_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n716_), .B2(new_n418_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n418_), .A2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n720_), .B2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n716_), .B2(new_n409_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n409_), .A2(G78gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n720_), .B2(new_n734_), .ZN(G1335gat));
  NOR3_X1   g534(.A1(new_n614_), .A2(new_n549_), .A3(new_n586_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n718_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n486_), .A3(new_n369_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n614_), .A2(new_n459_), .A3(new_n586_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n683_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n369_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n742_), .B2(new_n486_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n738_), .B2(new_n323_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n488_), .A2(new_n489_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n695_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n741_), .B2(new_n746_), .ZN(G1337gat));
  NAND2_X1  g546(.A1(new_n741_), .A2(new_n417_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n492_), .A2(new_n494_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n264_), .A2(new_n749_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n748_), .A2(G99gat), .B1(new_n738_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n493_), .A3(new_n393_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n683_), .A2(new_n393_), .A3(new_n740_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G106gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G106gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  NOR4_X1   g562(.A1(new_n264_), .A2(new_n323_), .A3(new_n412_), .A4(new_n393_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n719_), .A2(new_n765_), .A3(new_n460_), .A4(new_n614_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT54), .B1(new_n615_), .B2(new_n459_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n459_), .A2(new_n611_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n590_), .A2(new_n520_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n593_), .A2(new_n594_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(KEYINPUT55), .A3(new_n597_), .A4(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n587_), .A2(KEYINPUT12), .A3(new_n589_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT12), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n498_), .B2(new_n570_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n498_), .A2(new_n570_), .ZN(new_n776_));
  OAI22_X1  g575(.A1(new_n522_), .A2(new_n773_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n597_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT55), .B1(new_n595_), .B2(new_n597_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n608_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(new_n779_), .A3(new_n772_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n608_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n769_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n449_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n444_), .A2(new_n448_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n453_), .B2(new_n448_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n426_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI22_X1  g592(.A1(new_n451_), .A2(new_n454_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n609_), .A2(new_n611_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n549_), .B1(new_n789_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT57), .B(new_n549_), .C1(new_n789_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n793_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(new_n611_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n788_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n608_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n801_), .B(KEYINPUT58), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n798_), .B(new_n799_), .C1(new_n669_), .C2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n627_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n768_), .A2(KEYINPUT116), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT116), .B1(new_n768_), .B2(new_n810_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n764_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n813_), .A2(G113gat), .A3(new_n460_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n768_), .A2(new_n810_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n764_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n813_), .B2(KEYINPUT59), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n459_), .ZN(new_n820_));
  INV_X1    g619(.A(G113gat), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT117), .B(new_n815_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n819_), .B2(new_n459_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n814_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(new_n813_), .ZN(new_n827_));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n614_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(new_n829_), .C1(KEYINPUT60), .C2(new_n828_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n819_), .A2(new_n626_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g631(.A(G127gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n833_), .A3(new_n586_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n819_), .A2(new_n586_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n833_), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n827_), .A2(new_n837_), .A3(new_n624_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n819_), .A2(new_n670_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1343gat));
  OR2_X1    g639(.A1(new_n811_), .A2(new_n812_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n695_), .A2(new_n369_), .A3(new_n393_), .A4(new_n418_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT118), .Z(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n460_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT119), .B(G141gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1344gat));
  NOR2_X1   g646(.A1(new_n844_), .A2(new_n614_), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(G148gat), .Z(G1345gat));
  OAI21_X1  g648(.A(KEYINPUT120), .B1(new_n844_), .B2(new_n627_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n841_), .A2(new_n851_), .A3(new_n586_), .A4(new_n843_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n850_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1346gat));
  OAI21_X1  g655(.A(G162gat), .B1(new_n844_), .B2(new_n669_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n624_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n858_), .A2(G162gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n844_), .B2(new_n859_), .ZN(G1347gat));
  NOR3_X1   g659(.A1(new_n695_), .A2(new_n369_), .A3(new_n418_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n816_), .A2(new_n459_), .A3(new_n409_), .A4(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n286_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n202_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT122), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n868_), .A2(new_n869_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n866_), .A2(KEYINPUT122), .A3(new_n867_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n871_), .B2(new_n872_), .ZN(G1348gat));
  INV_X1    g672(.A(new_n816_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n861_), .A2(new_n409_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G176gat), .B1(new_n876_), .B2(new_n626_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n409_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT123), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n880_), .B(new_n409_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n861_), .A2(G176gat), .A3(new_n626_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n877_), .B1(new_n882_), .B2(new_n883_), .ZN(G1349gat));
  INV_X1    g683(.A(new_n280_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n885_), .A3(new_n586_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n861_), .A2(new_n586_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n879_), .B2(new_n881_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n886_), .B1(new_n888_), .B2(new_n213_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT124), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n891_), .B(new_n886_), .C1(new_n888_), .C2(new_n213_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1350gat));
  NAND4_X1  g692(.A1(new_n876_), .A2(new_n281_), .A3(new_n237_), .A4(new_n624_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n874_), .A2(new_n669_), .A3(new_n875_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n216_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n695_), .A2(new_n677_), .A3(new_n417_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n841_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n460_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n272_), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n614_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n273_), .ZN(G1353gat));
  INV_X1    g701(.A(new_n898_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n627_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT125), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n905_), .B(new_n907_), .ZN(G1354gat));
  AND3_X1   g707(.A1(new_n903_), .A2(G218gat), .A3(new_n670_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n898_), .A2(new_n858_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n910_), .A2(KEYINPUT126), .ZN(new_n911_));
  AOI21_X1  g710(.A(G218gat), .B1(new_n910_), .B2(KEYINPUT126), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n911_), .B2(new_n912_), .ZN(G1355gat));
endmodule


