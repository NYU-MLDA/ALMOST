//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT99), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT99), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT97), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  INV_X1    g009(.A(G197gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT97), .ZN(new_n212_));
  OAI21_X1  g011(.A(G204gat), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G211gat), .B(G218gat), .Z(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT21), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n208_), .A2(new_n213_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT100), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT100), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n208_), .A2(new_n213_), .A3(new_n221_), .A4(new_n218_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n215_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n211_), .A2(KEYINPUT97), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n209_), .A2(G197gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n203_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT98), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT99), .B(G204gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n211_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT98), .A4(new_n203_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n217_), .B1(new_n223_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  INV_X1    g036(.A(G141gat), .ZN(new_n238_));
  INV_X1    g037(.A(G148gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT95), .B1(new_n240_), .B2(KEYINPUT94), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(new_n240_), .B2(KEYINPUT95), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT96), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT2), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT2), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT96), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n246_), .A2(KEYINPUT96), .A3(G141gat), .A4(G148gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT95), .B(KEYINPUT3), .C1(new_n240_), .C2(KEYINPUT94), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259_));
  INV_X1    g058(.A(new_n255_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(KEYINPUT93), .A3(KEYINPUT1), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .A4(new_n254_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n240_), .A3(new_n248_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n237_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n234_), .A2(new_n236_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n215_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n211_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n203_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n221_), .B1(new_n272_), .B2(new_n218_), .ZN(new_n273_));
  NOR4_X1   g072(.A1(new_n270_), .A2(new_n271_), .A3(KEYINPUT100), .A4(KEYINPUT21), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n233_), .B(new_n269_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n216_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n258_), .A2(new_n266_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT29), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n235_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(G78gat), .B1(new_n268_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n236_), .B1(new_n234_), .B2(new_n267_), .ZN(new_n281_));
  INV_X1    g080(.A(G78gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n235_), .A3(new_n278_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n280_), .A2(G106gat), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(G106gat), .B1(new_n280_), .B2(new_n284_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n202_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G106gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n282_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n280_), .A2(new_n284_), .A3(G106gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT101), .A3(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n277_), .A2(KEYINPUT29), .ZN(new_n294_));
  INV_X1    g093(.A(G50gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT28), .B(G22gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(new_n293_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n300_), .A2(KEYINPUT101), .A3(new_n291_), .A4(new_n292_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT91), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n304_), .B(new_n305_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n303_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n241_), .A2(new_n242_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n256_), .B1(new_n309_), .B2(new_n252_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n265_), .A2(new_n240_), .A3(new_n248_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n258_), .A2(new_n307_), .A3(new_n266_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(KEYINPUT4), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n277_), .A2(new_n317_), .A3(new_n308_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT103), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n314_), .A2(KEYINPUT103), .A3(new_n316_), .A4(new_n318_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT104), .B(KEYINPUT0), .Z(new_n325_));
  XNOR2_X1  g124(.A(G1gat), .B(G29gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n321_), .A2(new_n329_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n334_));
  INV_X1    g133(.A(G190gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT87), .B1(new_n335_), .B2(KEYINPUT26), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT26), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(KEYINPUT26), .ZN(new_n341_));
  AND2_X1   g140(.A1(KEYINPUT86), .A2(G183gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(KEYINPUT86), .A2(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n340_), .B(new_n341_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT23), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n352_));
  AND2_X1   g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n351_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n346_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT86), .B(G183gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n344_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(KEYINPUT88), .A3(new_n340_), .A4(new_n341_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n349_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n358_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n351_), .B1(new_n362_), .B2(G190gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G169gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n334_), .B1(new_n276_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT25), .B(G183gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n338_), .A2(G190gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(new_n341_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n356_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n351_), .B1(G183gat), .B2(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n365_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n234_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n368_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT102), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n373_), .A2(KEYINPUT102), .A3(new_n365_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n372_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n334_), .B1(new_n276_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n378_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n234_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G64gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(G92gat), .Z(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(KEYINPUT32), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n378_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n381_), .A2(new_n382_), .B1(new_n356_), .B2(new_n371_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n378_), .B1(new_n234_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n368_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n333_), .A2(new_n394_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n393_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n399_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n386_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(new_n399_), .A3(new_n393_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n312_), .A2(KEYINPUT105), .A3(new_n313_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT105), .B1(new_n312_), .B2(new_n313_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n316_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n314_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n330_), .A3(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n406_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n332_), .B(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n402_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n302_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n404_), .A2(new_n405_), .A3(new_n403_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n393_), .B1(new_n379_), .B2(new_n388_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT27), .B1(new_n406_), .B2(new_n407_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n333_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n299_), .A3(new_n424_), .A4(new_n301_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G43gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT30), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(G71gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n361_), .A2(new_n432_), .A3(new_n366_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n361_), .B2(new_n366_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n367_), .A2(KEYINPUT89), .ZN(new_n436_));
  INV_X1    g235(.A(new_n431_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n361_), .A2(new_n432_), .A3(new_n366_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT90), .B(G99gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n435_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n428_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n435_), .A2(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n440_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n435_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n427_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n448_), .A3(KEYINPUT92), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT31), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT31), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n444_), .A2(new_n448_), .A3(KEYINPUT92), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n308_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n308_), .A3(new_n452_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n417_), .A2(new_n425_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n302_), .A2(new_n423_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT106), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n302_), .A2(KEYINPUT106), .A3(new_n423_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n455_), .A2(new_n424_), .A3(new_n456_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  INV_X1    g265(.A(G1gat), .ZN(new_n467_));
  INV_X1    g266(.A(G8gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT14), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G8gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G29gat), .ZN(new_n474_));
  INV_X1    g273(.A(G36gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G43gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G29gat), .A2(G36gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n477_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n480_), .A2(new_n295_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G43gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(G50gat), .B1(new_n484_), .B2(new_n479_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT74), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n295_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT74), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(G50gat), .A3(new_n479_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n486_), .A2(KEYINPUT15), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT15), .B1(new_n486_), .B2(new_n490_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n473_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT82), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n487_), .A2(KEYINPUT82), .A3(new_n489_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n472_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n493_), .A2(new_n494_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n497_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n473_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(KEYINPUT83), .A3(new_n498_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n494_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n504_), .A3(new_n473_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT84), .ZN(new_n509_));
  INV_X1    g308(.A(G169gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n211_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT85), .B1(new_n507_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n499_), .A2(new_n506_), .A3(new_n515_), .A4(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT64), .Z(new_n522_));
  INV_X1    g321(.A(KEYINPUT65), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n525_), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT67), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT6), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G99gat), .A3(G106gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT66), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(new_n539_), .A3(new_n530_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(G85gat), .A2(G92gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n529_), .A2(new_n537_), .A3(new_n530_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT8), .B1(new_n548_), .B2(new_n544_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT10), .B(G99gat), .Z(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n288_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n544_), .A2(KEYINPUT9), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n542_), .A2(new_n553_), .ZN(new_n554_));
  AND4_X1   g353(.A1(new_n537_), .A2(new_n551_), .A3(new_n552_), .A4(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT11), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n557_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n547_), .A2(new_n556_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT68), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n547_), .A2(new_n556_), .A3(KEYINPUT68), .A4(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n547_), .A2(new_n556_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n564_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n522_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n564_), .B(KEYINPUT70), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT69), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n547_), .A2(new_n556_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n572_), .A2(new_n576_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n566_), .A2(new_n522_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  NAND3_X1  g388(.A1(new_n574_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT72), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n573_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT72), .A3(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n594_), .A2(new_n589_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n465_), .A2(new_n520_), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n547_), .A2(new_n556_), .A3(new_n489_), .A4(new_n487_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT75), .ZN(new_n606_));
  OAI22_X1  g405(.A1(new_n579_), .A2(new_n580_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT76), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(KEYINPUT35), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT73), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n614_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n606_), .A2(new_n616_), .A3(new_n607_), .A4(new_n611_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(G134gat), .ZN(new_n620_));
  INV_X1    g419(.A(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n615_), .A2(new_n617_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n622_), .B(new_n618_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n615_), .A2(new_n625_), .A3(new_n617_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n627_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n626_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n472_), .B(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n575_), .B(KEYINPUT80), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G127gat), .B(G155gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(G183gat), .ZN(new_n641_));
  INV_X1    g440(.A(G211gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT17), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n638_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n636_), .A2(new_n565_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n636_), .A2(new_n565_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n647_), .A2(new_n645_), .A3(new_n648_), .A4(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n632_), .A2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT81), .Z(new_n654_));
  AND2_X1   g453(.A1(new_n604_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n467_), .A3(new_n333_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT38), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n462_), .A2(new_n464_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n457_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n624_), .A2(new_n626_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT107), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(KEYINPUT108), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n465_), .B2(new_n663_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n652_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n603_), .A2(new_n520_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n333_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n658_), .B1(new_n670_), .B2(G1gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n658_), .A3(G1gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n657_), .B1(new_n671_), .B2(new_n673_), .ZN(G1324gat));
  INV_X1    g473(.A(new_n423_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n655_), .A2(new_n468_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT39), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT108), .B1(new_n661_), .B2(new_n664_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n465_), .A2(new_n666_), .A3(new_n663_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n669_), .B(new_n651_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n677_), .B(G8gat), .C1(new_n680_), .C2(new_n423_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n668_), .A2(new_n669_), .A3(new_n675_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n677_), .B1(new_n683_), .B2(G8gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n676_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT40), .B(new_n676_), .C1(new_n682_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n456_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n308_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n655_), .A2(new_n690_), .A3(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n668_), .A2(new_n669_), .A3(new_n693_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT41), .B1(new_n695_), .B2(G15gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n302_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n655_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n668_), .A2(new_n669_), .A3(new_n701_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(G22gat), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n703_), .B2(G22gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n706_), .B2(new_n707_), .ZN(G1327gat));
  NOR2_X1   g507(.A1(new_n630_), .A2(new_n623_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n651_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n604_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G29gat), .B1(new_n712_), .B2(new_n333_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n632_), .B(KEYINPUT110), .ZN(new_n714_));
  OAI21_X1  g513(.A(KEYINPUT43), .B1(new_n465_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n632_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT43), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT111), .B1(new_n465_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n463_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n720_), .B(new_n717_), .C1(new_n721_), .C2(new_n457_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n715_), .A2(new_n719_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n669_), .A2(new_n652_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(KEYINPUT44), .A3(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(G29gat), .A3(new_n333_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n725_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n713_), .B1(new_n727_), .B2(new_n730_), .ZN(G1328gat));
  NAND4_X1  g530(.A1(new_n604_), .A2(new_n475_), .A3(new_n675_), .A4(new_n710_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT45), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n423_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n726_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT46), .B(new_n733_), .C1(new_n735_), .C2(new_n475_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n475_), .B1(new_n734_), .B2(new_n726_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n733_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n737_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1329gat));
  NAND4_X1  g540(.A1(new_n730_), .A2(G43gat), .A3(new_n693_), .A4(new_n726_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n693_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n477_), .B1(new_n711_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT47), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n747_), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1330gat));
  AOI21_X1  g548(.A(G50gat), .B1(new_n712_), .B2(new_n701_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n730_), .A2(G50gat), .A3(new_n726_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n701_), .ZN(G1331gat));
  NAND2_X1  g551(.A1(new_n603_), .A2(new_n520_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n465_), .A2(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(new_n654_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G57gat), .B1(new_n755_), .B2(new_n333_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n668_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n333_), .A2(G57gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1332gat));
  INV_X1    g560(.A(G64gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n762_), .A3(new_n675_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n675_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(G64gat), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n764_), .B2(G64gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n755_), .A2(new_n430_), .A3(new_n693_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G71gat), .B1(new_n758_), .B2(new_n743_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT49), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n771_), .A2(KEYINPUT49), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1334gat));
  NOR2_X1   g574(.A1(new_n302_), .A2(G78gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT112), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n755_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G78gat), .B1(new_n758_), .B2(new_n302_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(G1335gat));
  AND2_X1   g582(.A1(new_n754_), .A2(new_n710_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n333_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n753_), .A2(new_n651_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n723_), .A2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n424_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n790_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g590(.A(G92gat), .B1(new_n784_), .B2(new_n675_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n423_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n787_), .B2(new_n743_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n784_), .A2(new_n550_), .A3(new_n693_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g597(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n723_), .A2(new_n701_), .A3(new_n786_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G106gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT52), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n803_), .A3(G106gat), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n784_), .A2(new_n288_), .A3(new_n701_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n800_), .A2(new_n803_), .A3(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n800_), .B2(G106gat), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n799_), .B(new_n806_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n807_), .A2(new_n811_), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  NOR2_X1   g612(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n502_), .A2(new_n494_), .A3(new_n505_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n513_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT116), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n493_), .A2(new_n503_), .A3(new_n498_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n819_), .A3(new_n513_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n517_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n581_), .A2(new_n570_), .A3(new_n582_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n522_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n584_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n581_), .A2(new_n582_), .A3(KEYINPUT55), .A4(new_n583_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n589_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT72), .B1(new_n594_), .B2(new_n589_), .ZN(new_n835_));
  NOR4_X1   g634(.A1(new_n593_), .A2(new_n573_), .A3(new_n591_), .A4(new_n831_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n519_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n833_), .A3(KEYINPUT56), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n823_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n814_), .B1(new_n840_), .B2(new_n662_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n832_), .A2(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(new_n822_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n830_), .A2(new_n844_), .A3(new_n831_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n842_), .A2(new_n843_), .A3(new_n596_), .A4(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT118), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n596_), .A2(new_n845_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n822_), .B1(new_n832_), .B2(KEYINPUT56), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(new_n850_), .A3(KEYINPUT58), .A4(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n846_), .A2(new_n847_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n632_), .A4(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n814_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n839_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n856_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n709_), .B(new_n855_), .C1(new_n857_), .C2(new_n823_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n841_), .A2(new_n854_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n652_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n653_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n520_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT54), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n603_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n864_), .A2(new_n653_), .A3(new_n865_), .A4(new_n520_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n860_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n462_), .A2(new_n333_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n868_), .A2(new_n519_), .A3(new_n693_), .A4(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n520_), .A2(new_n873_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n868_), .A2(new_n693_), .A3(new_n870_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n859_), .A2(new_n652_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(new_n743_), .A3(new_n869_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n878_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n813_), .B1(new_n876_), .B2(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n880_), .A2(new_n881_), .A3(new_n879_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT59), .B1(new_n884_), .B2(KEYINPUT120), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n877_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n883_), .A2(new_n520_), .A3(new_n743_), .A4(new_n869_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT119), .B1(new_n891_), .B2(G113gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(KEYINPUT121), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n887_), .A2(new_n895_), .ZN(G1340gat));
  INV_X1    g695(.A(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n864_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n884_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n897_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n864_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n897_), .ZN(G1341gat));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n880_), .B2(new_n652_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT122), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n902_), .C1(new_n880_), .C2(new_n652_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n652_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(G127gat), .B2(new_n908_), .ZN(G1342gat));
  INV_X1    g708(.A(G134gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(new_n880_), .B2(new_n664_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT123), .B(new_n910_), .C1(new_n880_), .C2(new_n664_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n716_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(G134gat), .B2(new_n916_), .ZN(G1343gat));
  NOR3_X1   g716(.A1(new_n883_), .A2(new_n302_), .A3(new_n693_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(new_n333_), .A3(new_n423_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n520_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n238_), .ZN(G1344gat));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n864_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n239_), .ZN(G1345gat));
  INV_X1    g722(.A(new_n919_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n651_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT61), .B(G155gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1346gat));
  NOR3_X1   g726(.A1(new_n919_), .A2(new_n621_), .A3(new_n714_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n924_), .A2(new_n663_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n621_), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n423_), .A2(new_n333_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n883_), .A2(new_n743_), .A3(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT22), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n519_), .A4(new_n302_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(G169gat), .ZN(new_n937_));
  INV_X1    g736(.A(new_n933_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n938_), .A2(new_n520_), .A3(new_n701_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n510_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n937_), .B1(new_n941_), .B2(new_n936_), .ZN(G1348gat));
  NOR2_X1   g741(.A1(new_n938_), .A2(new_n701_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n603_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n933_), .A2(new_n302_), .A3(new_n651_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n362_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n933_), .A2(new_n302_), .A3(new_n369_), .A4(new_n651_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n947_), .B2(new_n949_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1350gat));
  NAND4_X1  g751(.A1(new_n943_), .A2(new_n370_), .A3(new_n341_), .A4(new_n663_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n933_), .A2(new_n302_), .A3(new_n632_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n954_), .A2(new_n955_), .A3(G190gat), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n954_), .B2(G190gat), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n953_), .B1(new_n956_), .B2(new_n957_), .ZN(G1351gat));
  AND2_X1   g757(.A1(new_n918_), .A2(new_n931_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n519_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n603_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(G204gat), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(new_n229_), .B2(new_n962_), .ZN(G1353gat));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n651_), .B1(new_n965_), .B2(new_n642_), .ZN(new_n966_));
  OR2_X1    g765(.A1(new_n966_), .A2(KEYINPUT126), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(KEYINPUT126), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n959_), .A2(new_n967_), .A3(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n965_), .A2(new_n642_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n969_), .B(new_n970_), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n918_), .A2(new_n663_), .A3(new_n931_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(G218gat), .ZN(new_n975_));
  NAND4_X1  g774(.A1(new_n918_), .A2(KEYINPUT127), .A3(new_n663_), .A4(new_n931_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n974_), .A2(new_n975_), .A3(new_n976_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n959_), .A2(G218gat), .A3(new_n632_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1355gat));
endmodule


