//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202_));
  XOR2_X1   g001(.A(G190gat), .B(G218gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G85gat), .B(G92gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n213_), .A2(new_n214_), .A3(new_n218_), .A4(new_n221_), .ZN(new_n222_));
  OAI22_X1  g021(.A1(new_n210_), .A2(new_n219_), .B1(new_n215_), .B2(G106gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT64), .B1(new_n223_), .B2(new_n212_), .ZN(new_n224_));
  OR4_X1    g023(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n217_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT7), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n209_), .A2(new_n225_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n220_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT8), .B1(new_n220_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n230_), .B2(new_n220_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n222_), .B(new_n224_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G29gat), .B(G36gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G43gat), .B(G50gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n237_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n245_), .A2(KEYINPUT72), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n237_), .A2(KEYINPUT67), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n231_), .B(new_n234_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n222_), .A2(new_n224_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n244_), .B(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n257_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n248_), .A2(new_n250_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n263_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n207_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n205_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(KEYINPUT36), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n268_), .A2(new_n271_), .A3(new_n264_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G15gat), .B(G22gat), .ZN(new_n279_));
  INV_X1    g078(.A(G1gat), .ZN(new_n280_));
  INV_X1    g079(.A(G8gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT14), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G8gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G231gat), .A2(G233gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n289_));
  XOR2_X1   g088(.A(G71gat), .B(G78gat), .Z(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n287_), .B(new_n296_), .Z(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT16), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT74), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G183gat), .B(G211gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT76), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n302_), .A2(KEYINPUT17), .ZN(new_n306_));
  INV_X1    g105(.A(new_n294_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n287_), .B(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(KEYINPUT17), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n202_), .B1(new_n278_), .B2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n253_), .A2(new_n257_), .A3(KEYINPUT12), .A4(new_n296_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT12), .B1(new_n237_), .B2(new_n307_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n237_), .A2(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G230gat), .A2(G233gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n237_), .B(new_n307_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n317_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G120gat), .B(G148gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT5), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G176gat), .B(G204gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT69), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI211_X1 g129(.A(KEYINPUT69), .B(new_n326_), .C1(new_n318_), .C2(new_n321_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n330_), .A2(KEYINPUT13), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT13), .B1(new_n330_), .B2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n311_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n276_), .A2(KEYINPUT77), .A3(new_n336_), .A4(new_n277_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n312_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n285_), .B(new_n244_), .Z(new_n341_));
  NAND2_X1  g140(.A1(G229gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n259_), .A2(new_n285_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT79), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(KEYINPUT79), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n285_), .A2(new_n244_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n349_), .B2(new_n342_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G141gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G169gat), .B(G197gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n312_), .A2(KEYINPUT78), .A3(new_n335_), .A4(new_n337_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n340_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT99), .ZN(new_n357_));
  AND2_X1   g156(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G169gat), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n360_), .A2(new_n361_), .B1(G169gat), .B2(G176gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT81), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT23), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n364_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n367_), .A2(KEYINPUT23), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT24), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(G169gat), .B2(G176gat), .ZN(new_n380_));
  OR2_X1    g179(.A1(G169gat), .A2(G176gat), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n378_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT26), .B(G190gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT25), .B(G183gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n377_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n374_), .A2(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT21), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(KEYINPUT21), .A3(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(G218gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G211gat), .ZN(new_n395_));
  INV_X1    g194(.A(G211gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G218gat), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n395_), .A2(new_n397_), .A3(KEYINPUT87), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT87), .B1(new_n395_), .B2(new_n397_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n392_), .B(new_n393_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n393_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n397_), .A3(KEYINPUT87), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n387_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n363_), .B1(G183gat), .B2(G190gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(new_n371_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n362_), .B1(new_n409_), .B2(new_n369_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(KEYINPUT25), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(KEYINPUT25), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n383_), .A3(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n414_), .A2(new_n382_), .A3(new_n368_), .A4(new_n372_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n410_), .A2(new_n415_), .A3(new_n400_), .A4(new_n404_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n406_), .A2(new_n416_), .A3(KEYINPUT20), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT19), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n410_), .A2(new_n415_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n405_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n419_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n374_), .A2(new_n400_), .A3(new_n386_), .A4(new_n404_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n420_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT27), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n417_), .A2(new_n419_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n424_), .A2(KEYINPUT20), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT96), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT96), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n424_), .A2(new_n439_), .A3(KEYINPUT20), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n422_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n436_), .B1(new_n441_), .B2(new_n419_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n435_), .B(KEYINPUT27), .C1(new_n430_), .C2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G141gat), .A2(G148gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT2), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(G141gat), .B2(G148gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G141gat), .A2(G148gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(KEYINPUT2), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n446_), .B(new_n449_), .C1(new_n451_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G155gat), .ZN(new_n455_));
  INV_X1    g254(.A(G162gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT83), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(G155gat), .B2(G162gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n457_), .B(new_n459_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(G141gat), .B(G148gat), .Z(new_n465_));
  AOI22_X1  g264(.A1(new_n454_), .A2(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT29), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT28), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT28), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G22gat), .B(G50gat), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n472_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n476_), .A2(G228gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(G228gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n405_), .A2(KEYINPUT85), .B1(G233gat), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n405_), .B1(new_n467_), .B2(new_n466_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G78gat), .B(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n475_), .B1(KEYINPUT88), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n483_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n485_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n486_), .B(new_n490_), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n445_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n421_), .B(KEYINPUT30), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G71gat), .B(G99gat), .ZN(new_n494_));
  INV_X1    g293(.A(G43gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G227gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(G15gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n493_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT31), .ZN(new_n502_));
  XOR2_X1   g301(.A(G127gat), .B(G134gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(G113gat), .B(G120gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  OR2_X1    g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT92), .B(G85gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G29gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT0), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n510_), .A2(KEYINPUT0), .ZN(new_n513_));
  OAI21_X1  g312(.A(G57gat), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n510_), .A2(KEYINPUT0), .ZN(new_n515_));
  INV_X1    g314(.A(G57gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(new_n511_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n509_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n517_), .A3(new_n509_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n505_), .A2(KEYINPUT4), .ZN(new_n523_));
  INV_X1    g322(.A(new_n466_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n503_), .B(new_n504_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n466_), .A2(new_n527_), .A3(KEYINPUT90), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n466_), .B2(KEYINPUT90), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT4), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT91), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n454_), .A2(new_n461_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n464_), .A2(new_n465_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT90), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n505_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n528_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT4), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n526_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n522_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n521_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n537_), .B2(KEYINPUT4), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT4), .ZN(new_n545_));
  AOI211_X1 g344(.A(KEYINPUT91), .B(new_n545_), .C1(new_n536_), .C2(new_n528_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n525_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n520_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(new_n518_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n541_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n492_), .A2(new_n508_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT98), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n491_), .A2(new_n551_), .A3(new_n444_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n547_), .A2(KEYINPUT33), .A3(new_n541_), .A4(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n522_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n522_), .B1(new_n536_), .B2(new_n528_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n549_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n556_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT94), .B1(new_n562_), .B2(new_n521_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n555_), .A2(new_n564_), .A3(new_n433_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT33), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n550_), .A2(KEYINPUT93), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT93), .B1(new_n550_), .B2(new_n566_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT95), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n565_), .B(new_n571_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n442_), .A2(KEYINPUT97), .A3(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n420_), .A2(new_n573_), .A3(new_n425_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT97), .B1(new_n442_), .B2(new_n573_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n551_), .A2(new_n574_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n554_), .B1(new_n578_), .B2(new_n491_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n508_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n553_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n491_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n555_), .A2(new_n564_), .A3(new_n433_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n550_), .A2(new_n566_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n550_), .A2(KEYINPUT93), .A3(new_n566_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n583_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n551_), .A2(new_n575_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n574_), .A2(new_n576_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n588_), .A2(new_n571_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n582_), .B1(new_n591_), .B2(new_n570_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT98), .B(new_n508_), .C1(new_n592_), .C2(new_n554_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n552_), .B1(new_n581_), .B2(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n356_), .A2(new_n357_), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n357_), .B1(new_n356_), .B2(new_n594_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n595_), .A2(new_n280_), .A3(new_n596_), .A4(new_n551_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT38), .ZN(new_n598_));
  INV_X1    g397(.A(new_n552_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n572_), .A2(new_n577_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n586_), .A2(new_n587_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n571_), .B1(new_n601_), .B2(new_n565_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n491_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n554_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT98), .B1(new_n605_), .B2(new_n508_), .ZN(new_n606_));
  AOI211_X1 g405(.A(new_n553_), .B(new_n580_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n599_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n273_), .B(KEYINPUT101), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n332_), .A2(new_n333_), .A3(new_n354_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT100), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n611_), .A2(new_n311_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n551_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n598_), .A2(new_n618_), .ZN(G1324gat));
  NOR2_X1   g418(.A1(new_n445_), .A2(G8gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n595_), .A2(new_n596_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n595_), .A2(KEYINPUT102), .A3(new_n596_), .A4(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n281_), .B1(new_n615_), .B2(new_n444_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n625_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1325gat));
  AOI21_X1  g431(.A(new_n498_), .B1(new_n615_), .B2(new_n580_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n634_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n595_), .A2(new_n498_), .A3(new_n596_), .A4(new_n580_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n615_), .B2(new_n582_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT42), .Z(new_n641_));
  NAND4_X1  g440(.A1(new_n595_), .A2(new_n639_), .A3(new_n596_), .A4(new_n582_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(new_n273_), .ZN(new_n644_));
  NOR4_X1   g443(.A1(new_n594_), .A2(new_n644_), .A3(new_n336_), .A4(new_n612_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n551_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT104), .B1(new_n614_), .B2(new_n336_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n613_), .A2(new_n648_), .A3(new_n311_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n278_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT105), .B(KEYINPUT43), .C1(new_n594_), .C2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n608_), .A2(new_n278_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT43), .B1(new_n655_), .B2(KEYINPUT105), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n651_), .B(KEYINPUT44), .C1(new_n654_), .C2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(G29gat), .A3(new_n551_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n654_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n650_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n646_), .B1(new_n658_), .B2(new_n661_), .ZN(G1328gat));
  XOR2_X1   g461(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n663_));
  INV_X1    g462(.A(G36gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n655_), .A2(KEYINPUT105), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n650_), .B1(new_n667_), .B2(new_n653_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n445_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n664_), .B1(new_n669_), .B2(new_n661_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n444_), .B(KEYINPUT106), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n645_), .A2(new_n664_), .A3(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT45), .Z(new_n674_));
  OAI21_X1  g473(.A(new_n663_), .B1(new_n670_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n657_), .A2(new_n444_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n668_), .A2(KEYINPUT44), .ZN(new_n677_));
  OAI21_X1  g476(.A(G36gat), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n674_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n663_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n681_), .ZN(G1329gat));
  NAND2_X1  g481(.A1(new_n645_), .A2(new_n580_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(new_n495_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n657_), .A2(G43gat), .A3(new_n580_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n677_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT47), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n688_), .B(new_n684_), .C1(new_n685_), .C2(new_n677_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1330gat));
  INV_X1    g489(.A(G50gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n645_), .A2(new_n691_), .A3(new_n582_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n491_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n661_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G50gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n693_), .B2(new_n661_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n692_), .B1(new_n696_), .B2(new_n697_), .ZN(G1331gat));
  NOR3_X1   g497(.A1(new_n594_), .A2(new_n354_), .A3(new_n335_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(new_n312_), .A3(new_n337_), .ZN(new_n700_));
  AOI211_X1 g499(.A(KEYINPUT109), .B(G57gat), .C1(new_n700_), .C2(new_n551_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n551_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n516_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n354_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n336_), .A2(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n611_), .A2(new_n335_), .A3(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n617_), .A2(new_n516_), .ZN(new_n708_));
  AOI211_X1 g507(.A(new_n701_), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n707_), .B2(new_n672_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT48), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n700_), .A2(new_n710_), .A3(new_n672_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n707_), .B2(new_n580_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT49), .Z(new_n717_));
  NOR2_X1   g516(.A1(new_n508_), .A2(G71gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT110), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n700_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1334gat));
  INV_X1    g520(.A(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n707_), .B2(new_n582_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n700_), .A2(new_n722_), .A3(new_n582_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1335gat));
  AND3_X1   g525(.A1(new_n699_), .A2(new_n273_), .A3(new_n311_), .ZN(new_n727_));
  INV_X1    g526(.A(G85gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n551_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n335_), .A2(new_n336_), .A3(new_n354_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n656_), .B2(new_n654_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT111), .B(new_n730_), .C1(new_n656_), .C2(new_n654_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n617_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n729_), .B1(new_n735_), .B2(new_n728_), .ZN(G1336gat));
  INV_X1    g535(.A(G92gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n727_), .A2(new_n737_), .A3(new_n444_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n671_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n737_), .ZN(G1337gat));
  NAND3_X1  g539(.A1(new_n727_), .A2(new_n580_), .A3(new_n216_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n508_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n227_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT51), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n745_), .B(new_n741_), .C1(new_n742_), .C2(new_n227_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n727_), .A2(new_n217_), .A3(new_n582_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n582_), .B(new_n730_), .C1(new_n656_), .C2(new_n654_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G106gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G106gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT53), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n748_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1339gat));
  NOR3_X1   g556(.A1(new_n492_), .A2(new_n508_), .A3(new_n617_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n330_), .A2(new_n331_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n350_), .A2(new_n353_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n349_), .A2(new_n342_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n353_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT117), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n760_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767_));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n318_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n318_), .B2(new_n768_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n313_), .A2(new_n316_), .A3(KEYINPUT55), .A4(new_n317_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n313_), .A2(new_n316_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n320_), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT114), .B(new_n317_), .C1(new_n313_), .C2(new_n316_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT115), .B(new_n325_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n354_), .A2(new_n327_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n772_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n774_), .A2(new_n320_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT114), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n774_), .A2(new_n773_), .A3(new_n320_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n318_), .A2(new_n768_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT113), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n318_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n326_), .B1(new_n787_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT115), .B1(new_n793_), .B2(KEYINPUT116), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n782_), .B1(new_n792_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n766_), .B1(new_n780_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n797_), .B2(new_n644_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n765_), .A2(new_n327_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n793_), .B(new_n325_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n325_), .B1(new_n771_), .B2(new_n777_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n803_), .A4(new_n801_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n278_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n644_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n799_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n798_), .A2(KEYINPUT118), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n311_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n652_), .A2(new_n335_), .A3(new_n336_), .A4(new_n705_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n759_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  INV_X1    g618(.A(new_n817_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n808_), .A2(new_n278_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n765_), .A2(new_n327_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n806_), .B2(KEYINPUT56), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT58), .B1(new_n824_), .B2(new_n803_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n821_), .B1(new_n798_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n781_), .B1(new_n806_), .B2(new_n794_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT116), .B1(new_n792_), .B2(KEYINPUT115), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(KEYINPUT56), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n273_), .B1(new_n830_), .B2(new_n766_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n809_), .B(KEYINPUT119), .C1(new_n831_), .C2(KEYINPUT57), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(new_n832_), .A3(new_n810_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n820_), .B1(new_n833_), .B2(new_n311_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n759_), .A2(KEYINPUT59), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n818_), .A2(new_n819_), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n705_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n810_), .A2(new_n809_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n840_), .B(KEYINPUT57), .C1(new_n797_), .C2(new_n644_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n812_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n336_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n758_), .B1(new_n844_), .B2(new_n820_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n705_), .A2(G113gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n838_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n833_), .A2(new_n311_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n817_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n845_), .A2(KEYINPUT59), .B1(new_n851_), .B2(new_n835_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n852_), .B2(new_n334_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n334_), .A2(new_n854_), .A3(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n854_), .B2(new_n849_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n818_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n848_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G120gat), .B1(new_n837_), .B2(new_n335_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n852_), .B2(new_n336_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n845_), .A2(G127gat), .A3(new_n311_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT121), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G127gat), .B1(new_n837_), .B2(new_n311_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  INV_X1    g667(.A(new_n865_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n870_), .ZN(G1342gat));
  OAI21_X1  g670(.A(G134gat), .B1(new_n837_), .B2(new_n652_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n610_), .A2(G134gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n845_), .B2(new_n873_), .ZN(G1343gat));
  NAND2_X1  g673(.A1(new_n813_), .A2(new_n817_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n580_), .A2(new_n491_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n672_), .A2(new_n617_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n879_), .A2(G141gat), .A3(new_n705_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G141gat), .B1(new_n879_), .B2(new_n705_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1344gat));
  XOR2_X1   g681(.A(KEYINPUT122), .B(G148gat), .Z(new_n883_));
  OR3_X1    g682(.A1(new_n879_), .A2(new_n335_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n879_), .B2(new_n335_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1345gat));
  NAND3_X1  g685(.A1(new_n877_), .A2(new_n336_), .A3(new_n878_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n879_), .B2(new_n652_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n609_), .A2(new_n456_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n879_), .B2(new_n891_), .ZN(G1347gat));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n671_), .A2(new_n551_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n580_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n582_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n851_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n705_), .ZN(new_n898_));
  INV_X1    g697(.A(G169gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n893_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT62), .B(G169gat), .C1(new_n897_), .C2(new_n705_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n361_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  INV_X1    g702(.A(new_n897_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n334_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n582_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n334_), .A2(G176gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n895_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n905_), .A2(new_n360_), .B1(new_n906_), .B2(new_n908_), .ZN(G1349gat));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n895_), .A2(new_n311_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n906_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(G183gat), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n311_), .A2(new_n384_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n897_), .A2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n910_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  OAI221_X1 g715(.A(KEYINPUT123), .B1(new_n897_), .B2(new_n914_), .C1(new_n912_), .C2(G183gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n897_), .B2(new_n652_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n904_), .A2(new_n383_), .A3(new_n609_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1351gat));
  NAND3_X1  g722(.A1(new_n877_), .A2(new_n354_), .A3(new_n894_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n875_), .A2(new_n334_), .A3(new_n876_), .A4(new_n894_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n927_), .A2(new_n928_), .A3(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n928_), .B1(new_n927_), .B2(new_n930_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n926_), .B1(new_n932_), .B2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n927_), .A2(new_n930_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(KEYINPUT126), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n936_), .A2(KEYINPUT125), .A3(G204gat), .A4(new_n931_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(G1353gat));
  AND3_X1   g737(.A1(new_n877_), .A2(new_n336_), .A3(new_n894_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  AND2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n939_), .B2(new_n940_), .ZN(G1354gat));
  AND2_X1   g742(.A1(new_n877_), .A2(new_n894_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n609_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n278_), .A2(G218gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT127), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n945_), .A2(new_n394_), .B1(new_n944_), .B2(new_n947_), .ZN(G1355gat));
endmodule


