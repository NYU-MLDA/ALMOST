//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT86), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT22), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G169gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT86), .A2(G176gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT84), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT84), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n219_), .B2(KEYINPUT23), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n218_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n216_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n229_));
  AND2_X1   g028(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n231_));
  OAI22_X1  g030(.A1(new_n228_), .A2(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n206_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(KEYINPUT98), .A2(KEYINPUT24), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT98), .A2(KEYINPUT24), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n234_), .B(new_n235_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT99), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n232_), .A2(new_n238_), .A3(KEYINPUT99), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n244_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n227_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G218gat), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n247_), .A2(G211gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(G211gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT21), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT96), .B(G204gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G197gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT95), .B(G197gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G204gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n250_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n248_), .A2(new_n249_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  OAI22_X1  g056(.A1(G197gat), .A2(new_n251_), .B1(new_n253_), .B2(G204gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT21), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n255_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n204_), .B1(new_n246_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT101), .ZN(new_n264_));
  OAI21_X1  g063(.A(G169gat), .B1(new_n208_), .B2(KEYINPUT85), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n206_), .A3(KEYINPUT22), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n265_), .A2(new_n267_), .A3(new_n205_), .A4(new_n210_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n215_), .ZN(new_n269_));
  AND2_X1   g068(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT82), .B(G190gat), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n272_), .A2(new_n273_), .B1(new_n220_), .B2(new_n218_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  OR3_X1    g074(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n235_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n212_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n228_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n273_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n231_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT25), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n272_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n275_), .B1(new_n288_), .B2(new_n224_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n264_), .B1(new_n289_), .B2(new_n262_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n263_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n253_), .A2(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(G204gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT96), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT96), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G204gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(G197gat), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT21), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n261_), .A3(new_n256_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n255_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n287_), .A2(new_n284_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n276_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n280_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n215_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n224_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n272_), .A2(new_n273_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n220_), .A2(new_n218_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n268_), .A3(new_n215_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n301_), .A2(new_n311_), .A3(KEYINPUT101), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n203_), .B1(new_n291_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT20), .B1(new_n301_), .B2(new_n311_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n203_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT100), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n246_), .A2(new_n262_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n242_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT99), .B1(new_n232_), .B2(new_n238_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n245_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n224_), .A2(new_n226_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n216_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT100), .B1(new_n326_), .B2(new_n301_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n316_), .B(new_n317_), .C1(new_n319_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n314_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT18), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n316_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n203_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n322_), .A2(new_n325_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT20), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT101), .B1(new_n301_), .B2(new_n311_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT102), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n317_), .A4(new_n312_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n263_), .A2(new_n290_), .A3(new_n317_), .A4(new_n312_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT102), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n338_), .A2(new_n344_), .A3(new_n346_), .A4(new_n334_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n336_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n349_));
  INV_X1    g148(.A(G155gat), .ZN(new_n350_));
  INV_X1    g149(.A(G162gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT1), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(G155gat), .A3(G162gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT91), .B1(G155gat), .B2(G162gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n352_), .A2(new_n354_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G141gat), .B(G148gat), .Z(new_n359_));
  AND3_X1   g158(.A1(new_n358_), .A2(KEYINPUT92), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT92), .B1(new_n358_), .B2(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n352_), .A2(new_n357_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n353_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n365_));
  INV_X1    g164(.A(G141gat), .ZN(new_n366_));
  INV_X1    g165(.A(G148gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT3), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n365_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n368_), .A2(new_n370_), .ZN(new_n377_));
  AND3_X1   g176(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n372_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n379_), .A3(KEYINPUT93), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n364_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT94), .B1(new_n362_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n361_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n358_), .A2(KEYINPUT92), .A3(new_n359_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n377_), .A2(new_n379_), .A3(KEYINPUT93), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT93), .B1(new_n377_), .B2(new_n379_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n363_), .B(new_n353_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G127gat), .B(G134gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n382_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  OR3_X1    g193(.A1(new_n362_), .A2(new_n381_), .A3(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT103), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G85gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n394_), .A2(KEYINPUT4), .A3(new_n395_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n382_), .A2(new_n390_), .A3(new_n406_), .A4(new_n393_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n397_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n399_), .B(new_n404_), .C1(new_n405_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT104), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n399_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n403_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n394_), .A2(KEYINPUT4), .A3(new_n395_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(new_n397_), .A3(new_n407_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT104), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n399_), .A4(new_n404_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n410_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n348_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(new_n398_), .A3(new_n407_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n394_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n421_), .A2(new_n403_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n409_), .A2(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n338_), .A2(new_n344_), .A3(new_n346_), .A4(new_n333_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n333_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n318_), .B1(new_n246_), .B2(new_n262_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n326_), .A2(new_n301_), .A3(KEYINPUT100), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n315_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n317_), .A2(new_n428_), .B1(new_n345_), .B2(KEYINPUT102), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n345_), .A2(KEYINPUT102), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n425_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n414_), .A2(KEYINPUT33), .A3(new_n399_), .A4(new_n404_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n423_), .A2(new_n424_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n418_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G22gat), .B(G50gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n382_), .A2(new_n390_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT28), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n435_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n435_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n439_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G78gat), .B(G106gat), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n382_), .A2(new_n390_), .A3(KEYINPUT29), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n262_), .B1(G228gat), .B2(G233gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT97), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n453_), .A3(new_n450_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n438_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n456_));
  OAI211_X1 g255(.A(G228gat), .B(G233gat), .C1(new_n456_), .C2(new_n262_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n448_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n449_), .A2(new_n453_), .A3(new_n450_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n453_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n448_), .B(new_n457_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n446_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n447_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(new_n445_), .A3(new_n442_), .A4(new_n461_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n434_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n417_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n431_), .A2(new_n424_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n329_), .B2(new_n425_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n471_), .A2(new_n472_), .B1(new_n424_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n311_), .B(KEYINPUT30), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G71gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G99gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(G15gat), .B(G43gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT87), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n483_), .B(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n480_), .A3(new_n486_), .ZN(new_n487_));
  OR3_X1    g286(.A1(new_n477_), .A2(new_n486_), .A3(new_n478_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n393_), .B(KEYINPUT31), .Z(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT89), .Z(new_n491_));
  NAND4_X1  g290(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT90), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n490_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n492_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n474_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(new_n467_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n496_), .A2(new_n417_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n476_), .A2(new_n496_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(G190gat), .B(G218gat), .Z(new_n501_));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT36), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT65), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT65), .B1(new_n508_), .B2(new_n510_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI221_X1 g312(.A(KEYINPUT66), .B1(KEYINPUT67), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT66), .B1(KEYINPUT67), .B2(KEYINPUT7), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n514_), .B(new_n517_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n506_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n515_), .A2(new_n516_), .B1(KEYINPUT66), .B2(KEYINPUT7), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n515_), .A2(new_n516_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(KEYINPUT68), .C1(new_n511_), .C2(new_n512_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G85gat), .B(G92gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n519_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n519_), .A2(new_n523_), .A3(KEYINPUT69), .A4(new_n525_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n508_), .A2(new_n510_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT70), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n508_), .A2(new_n510_), .A3(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n522_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n524_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n528_), .A2(new_n529_), .A3(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G29gat), .B(G36gat), .Z(new_n540_));
  XOR2_X1   g339(.A(G43gat), .B(G50gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n513_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n536_), .A2(KEYINPUT9), .ZN(new_n544_));
  INV_X1    g343(.A(G85gat), .ZN(new_n545_));
  INV_X1    g344(.A(G92gat), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT9), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT10), .B(G99gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT64), .B(G106gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n543_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n539_), .A2(new_n542_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n554_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n542_), .B(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n539_), .B2(new_n551_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n557_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n560_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n551_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n537_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n529_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n555_), .B1(new_n568_), .B2(new_n542_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n539_), .A2(new_n551_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n565_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n505_), .B1(new_n564_), .B2(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n539_), .A2(new_n542_), .A3(new_n551_), .ZN(new_n575_));
  OAI211_X1 g374(.A(KEYINPUT35), .B(new_n554_), .C1(new_n575_), .C2(new_n563_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n565_), .A3(new_n572_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n503_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT75), .Z(new_n580_));
  NAND3_X1  g379(.A1(new_n576_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n500_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584_));
  INV_X1    g383(.A(G1gat), .ZN(new_n585_));
  INV_X1    g384(.A(G8gat), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT14), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G1gat), .B(G8gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n542_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT80), .Z(new_n595_));
  OR2_X1    g394(.A1(new_n562_), .A2(new_n590_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n542_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n602_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT73), .ZN(new_n606_));
  XOR2_X1   g405(.A(G57gat), .B(G64gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT71), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT11), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G71gat), .B(G78gat), .Z(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n609_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(new_n613_), .A3(new_n611_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n570_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n614_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n568_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(G230gat), .B(G233gat), .C1(new_n616_), .C2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n570_), .A2(new_n615_), .A3(KEYINPUT12), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n568_), .B2(new_n617_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n568_), .A2(new_n617_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n620_), .A2(new_n622_), .A3(new_n623_), .A4(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n619_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT5), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n628_), .B(new_n629_), .Z(new_n630_));
  OAI21_X1  g429(.A(new_n606_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n630_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n619_), .A2(new_n625_), .A3(KEYINPUT73), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n630_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(KEYINPUT13), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT13), .B1(new_n634_), .B2(new_n635_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n590_), .B(new_n639_), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n617_), .B(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(G127gat), .B(G155gat), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT16), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT17), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n641_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT17), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n641_), .A2(new_n648_), .A3(new_n645_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT78), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(KEYINPUT78), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n583_), .A2(new_n605_), .A3(new_n638_), .A4(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n417_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT105), .Z(new_n656_));
  INV_X1    g455(.A(new_n605_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n634_), .A2(new_n635_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT13), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n634_), .A2(KEYINPUT13), .A3(new_n635_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT76), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n576_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n504_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT77), .B1(new_n574_), .B2(new_n581_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT37), .B(new_n666_), .C1(new_n667_), .C2(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT77), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT37), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT76), .A3(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n652_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n662_), .A2(new_n673_), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n657_), .B(new_n500_), .C1(new_n674_), .C2(KEYINPUT79), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(KEYINPUT79), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n675_), .A2(new_n585_), .A3(new_n417_), .A4(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT38), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n656_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT106), .ZN(G1324gat));
  NAND4_X1  g479(.A1(new_n675_), .A2(new_n586_), .A3(new_n497_), .A4(new_n676_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT107), .ZN(new_n682_));
  OAI21_X1  g481(.A(G8gat), .B1(new_n653_), .B2(new_n474_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT39), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(G1325gat));
  OAI21_X1  g486(.A(G15gat), .B1(new_n653_), .B2(new_n496_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT41), .Z(new_n689_));
  NAND2_X1  g488(.A1(new_n675_), .A2(new_n676_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n496_), .A2(G15gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(G1326gat));
  XNOR2_X1  g491(.A(new_n467_), .B(KEYINPUT108), .ZN(new_n693_));
  OAI21_X1  g492(.A(G22gat), .B1(new_n653_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT42), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n693_), .A2(G22gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n690_), .B2(new_n696_), .ZN(G1327gat));
  NOR2_X1   g496(.A1(new_n500_), .A2(new_n657_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n582_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n652_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n638_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(G29gat), .A3(new_n654_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n652_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n638_), .A2(new_n605_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n663_), .B1(new_n582_), .B2(new_n669_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n666_), .A2(KEYINPUT37), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n672_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n668_), .A2(new_n712_), .A3(new_n672_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n499_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n434_), .A2(new_n468_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n496_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n707_), .B1(new_n714_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT43), .B1(new_n668_), .B2(new_n672_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n706_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n668_), .A2(new_n712_), .A3(new_n672_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n712_), .B1(new_n668_), .B2(new_n672_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n718_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT43), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n705_), .B1(new_n729_), .B2(new_n721_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n725_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n706_), .B1(new_n719_), .B2(new_n722_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n417_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n703_), .B1(new_n736_), .B2(G29gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT111), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n702_), .A2(G36gat), .A3(new_n474_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT45), .Z(new_n740_));
  AOI21_X1  g539(.A(new_n474_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT110), .B1(new_n730_), .B2(KEYINPUT44), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n728_), .A2(KEYINPUT43), .B1(new_n718_), .B2(new_n720_), .ZN(new_n743_));
  NOR4_X1   g542(.A1(new_n743_), .A2(new_n724_), .A3(new_n734_), .A4(new_n705_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n741_), .B(KEYINPUT112), .C1(new_n742_), .C2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G36gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT112), .B1(new_n732_), .B2(new_n741_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n740_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT46), .B(new_n740_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1329gat));
  AND4_X1   g551(.A1(G43gat), .A2(new_n732_), .A3(new_n717_), .A4(new_n735_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n755_));
  INV_X1    g554(.A(new_n702_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n717_), .ZN(new_n757_));
  INV_X1    g556(.A(G43gat), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n755_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n759_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT47), .B1(new_n753_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1330gat));
  INV_X1    g562(.A(new_n693_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G50gat), .B1(new_n756_), .B2(new_n764_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n732_), .A2(new_n735_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n467_), .A2(G50gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(G1331gat));
  NOR2_X1   g567(.A1(new_n704_), .A2(new_n605_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n583_), .A2(new_n662_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n583_), .A2(KEYINPUT113), .A3(new_n662_), .A4(new_n769_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G57gat), .B1(new_n654_), .B2(KEYINPUT114), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n774_), .B(new_n775_), .C1(KEYINPUT114), .C2(G57gat), .ZN(new_n776_));
  INV_X1    g575(.A(G57gat), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n500_), .A2(new_n605_), .A3(new_n638_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n673_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n654_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n776_), .A2(new_n781_), .ZN(G1332gat));
  OR3_X1    g581(.A1(new_n780_), .A2(G64gat), .A3(new_n474_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n772_), .A2(new_n497_), .A3(new_n773_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT48), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G64gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G64gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT115), .ZN(G1333gat));
  NAND2_X1  g588(.A1(new_n774_), .A2(new_n717_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G71gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT49), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n496_), .A2(G71gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n780_), .B2(new_n793_), .ZN(G1334gat));
  INV_X1    g593(.A(G78gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n774_), .B2(new_n764_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n764_), .A2(new_n795_), .ZN(new_n800_));
  OAI22_X1  g599(.A1(new_n798_), .A2(new_n799_), .B1(new_n780_), .B2(new_n800_), .ZN(G1335gat));
  NAND3_X1  g600(.A1(new_n662_), .A2(new_n657_), .A3(new_n704_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n743_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803_), .B2(new_n654_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n778_), .A2(new_n700_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n545_), .A3(new_n417_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(G1336gat));
  OAI21_X1  g607(.A(G92gat), .B1(new_n803_), .B2(new_n474_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n546_), .A3(new_n497_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n803_), .B2(new_n496_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n717_), .A2(new_n548_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n805_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n806_), .A2(new_n549_), .A3(new_n467_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G106gat), .B1(new_n803_), .B2(new_n468_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT53), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n816_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n674_), .B2(new_n657_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n662_), .A2(new_n673_), .A3(KEYINPUT117), .A4(new_n605_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n779_), .A2(new_n638_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT117), .B1(new_n830_), .B2(new_n605_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n674_), .A2(new_n826_), .A3(new_n657_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(KEYINPUT54), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n829_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n710_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n596_), .A2(new_n597_), .A3(new_n593_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n591_), .A2(new_n592_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n602_), .A3(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n603_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n634_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n625_), .A2(KEYINPUT118), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n625_), .B2(new_n842_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n625_), .A2(new_n842_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n620_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(G230gat), .A3(G233gat), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .A4(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n630_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n848_), .B2(new_n630_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n841_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n835_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT58), .B(new_n841_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n605_), .B(new_n634_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n658_), .A2(new_n839_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n582_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(KEYINPUT57), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(KEYINPUT57), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n704_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n834_), .A2(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n497_), .A2(new_n654_), .A3(new_n496_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(KEYINPUT59), .A3(new_n468_), .A4(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n634_), .A2(new_n605_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n848_), .A2(new_n630_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n630_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n857_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n699_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n866_), .A2(new_n874_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n652_), .B1(new_n875_), .B2(new_n860_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n829_), .A2(new_n833_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n468_), .B(new_n864_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n657_), .B1(new_n865_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(G113gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n605_), .A2(new_n882_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n881_), .A2(new_n882_), .B1(new_n878_), .B2(new_n883_), .ZN(G1340gat));
  AOI21_X1  g683(.A(new_n638_), .B1(new_n865_), .B2(new_n880_), .ZN(new_n885_));
  INV_X1    g684(.A(G120gat), .ZN(new_n886_));
  INV_X1    g685(.A(new_n878_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n888_));
  AOI21_X1  g687(.A(G120gat), .B1(new_n662_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n886_), .A2(KEYINPUT60), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(KEYINPUT119), .B1(new_n887_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  NOR4_X1   g692(.A1(new_n878_), .A2(new_n893_), .A3(new_n890_), .A4(new_n889_), .ZN(new_n894_));
  OAI22_X1  g693(.A1(new_n885_), .A2(new_n886_), .B1(new_n892_), .B2(new_n894_), .ZN(G1341gat));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n878_), .B2(new_n704_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT120), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n899_), .B(new_n896_), .C1(new_n878_), .C2(new_n704_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n865_), .A2(new_n880_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n704_), .A2(new_n896_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n898_), .A2(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1342gat));
  INV_X1    g702(.A(G134gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n887_), .A2(new_n904_), .A3(new_n582_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n835_), .B1(new_n865_), .B2(new_n880_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1343gat));
  NOR4_X1   g706(.A1(new_n497_), .A2(new_n717_), .A3(new_n468_), .A4(new_n654_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n834_), .B2(new_n862_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n605_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n662_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n652_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1346gat));
  NAND2_X1  g716(.A1(new_n910_), .A2(new_n582_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n351_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n351_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n910_), .A2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n920_), .A3(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n922_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G162gat), .B1(new_n910_), .B2(new_n582_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n926_), .ZN(G1347gat));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n499_), .A2(new_n497_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n764_), .A2(new_n929_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n605_), .B(new_n930_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n931_), .B2(G169gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n928_), .A3(G169gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(KEYINPUT62), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n207_), .A2(new_n209_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n931_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n932_), .A2(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n935_), .A2(new_n939_), .ZN(G1348gat));
  NAND3_X1  g739(.A1(new_n863_), .A2(new_n662_), .A3(new_n930_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n205_), .A2(new_n210_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(KEYINPUT123), .A3(new_n942_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n876_), .A2(new_n877_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n467_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n638_), .A2(new_n233_), .A3(new_n929_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n945_), .A2(new_n946_), .B1(new_n948_), .B2(new_n949_), .ZN(G1349gat));
  NAND4_X1  g749(.A1(new_n948_), .A2(new_n652_), .A3(new_n497_), .A4(new_n499_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n947_), .A2(new_n764_), .A3(new_n929_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n704_), .A2(new_n231_), .A3(new_n230_), .ZN(new_n953_));
  AOI22_X1  g752(.A1(new_n951_), .A2(new_n272_), .B1(new_n952_), .B2(new_n953_), .ZN(G1350gat));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n710_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(G190gat), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n582_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(KEYINPUT124), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n952_), .A2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n956_), .A2(new_n959_), .ZN(G1351gat));
  AND3_X1   g759(.A1(new_n497_), .A2(new_n470_), .A3(new_n496_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n863_), .A2(new_n605_), .A3(new_n961_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g762(.A1(new_n863_), .A2(new_n662_), .A3(new_n961_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n964_), .A2(new_n251_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n965_), .B1(new_n293_), .B2(new_n964_), .ZN(G1353gat));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n967_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968_));
  AOI211_X1 g767(.A(new_n968_), .B(new_n704_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n863_), .A2(new_n961_), .A3(new_n969_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n967_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n971_));
  XOR2_X1   g770(.A(new_n971_), .B(KEYINPUT126), .Z(new_n972_));
  XNOR2_X1  g771(.A(new_n970_), .B(new_n972_), .ZN(G1354gat));
  OAI211_X1 g772(.A(new_n582_), .B(new_n961_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n975_), .A2(G218gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n977_));
  AND2_X1   g776(.A1(new_n863_), .A2(new_n961_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n835_), .A2(new_n247_), .ZN(new_n979_));
  AOI22_X1  g778(.A1(new_n976_), .A2(new_n977_), .B1(new_n978_), .B2(new_n979_), .ZN(G1355gat));
endmodule


