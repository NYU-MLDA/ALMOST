//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n967_, new_n968_, new_n969_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT79), .B(G43gat), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT30), .ZN(new_n209_));
  NOR3_X1   g008(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(G169gat), .B2(G176gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT25), .B(G183gat), .Z(new_n218_));
  OAI21_X1  g017(.A(new_n215_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT23), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n220_), .A2(new_n222_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(KEYINPUT23), .A3(new_n226_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n209_), .B1(new_n229_), .B2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n231_), .A2(new_n232_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n238_), .B1(new_n242_), .B2(new_n230_), .ZN(new_n243_));
  OAI221_X1 g042(.A(new_n215_), .B1(new_n217_), .B2(new_n218_), .C1(new_n223_), .C2(new_n227_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(KEYINPUT30), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G99gat), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n241_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n241_), .B2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n208_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n229_), .A2(new_n240_), .A3(new_n209_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT30), .B1(new_n243_), .B2(new_n244_), .ZN(new_n251_));
  OAI21_X1  g050(.A(G99gat), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n241_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n207_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255_));
  INV_X1    g054(.A(G15gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G71gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT80), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n249_), .B2(new_n254_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n206_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G57gat), .B(G85gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT91), .ZN(new_n264_));
  INV_X1    g063(.A(G1gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT92), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G29gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n266_), .A2(new_n269_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n202_), .B(new_n203_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT3), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n276_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(KEYINPUT1), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(G155gat), .A3(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n289_), .A3(new_n283_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291_));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n273_), .B(new_n286_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n286_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n204_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n297_), .A3(KEYINPUT4), .ZN(new_n300_));
  INV_X1    g099(.A(new_n298_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n300_), .B(new_n301_), .C1(KEYINPUT4), .C2(new_n297_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n272_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n272_), .A2(new_n302_), .A3(new_n299_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n249_), .A2(new_n254_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n258_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(KEYINPUT80), .A3(new_n259_), .A4(new_n205_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n262_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT84), .B1(new_n312_), .B2(G197gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n314_));
  INV_X1    g113(.A(G197gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(G197gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT87), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n313_), .A2(new_n316_), .A3(new_n320_), .A4(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT21), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G218gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G211gat), .ZN(new_n327_));
  INV_X1    g126(.A(G211gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G218gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT86), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n322_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n316_), .A2(new_n317_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .A4(new_n313_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n313_), .A2(new_n316_), .A3(new_n336_), .A4(new_n317_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT85), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n315_), .A2(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n317_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n330_), .B1(KEYINPUT21), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n344_), .A2(KEYINPUT83), .B1(G228gat), .B2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n290_), .A2(new_n291_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT81), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n348_), .A2(new_n349_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n344_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n345_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(G22gat), .B(G50gat), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n346_), .A3(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n296_), .B2(KEYINPUT29), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n359_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n353_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n357_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n358_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n353_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT88), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n352_), .A2(new_n362_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n352_), .B1(new_n362_), .B2(new_n369_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT19), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n218_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT25), .B(G183gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT89), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n216_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n213_), .A2(new_n211_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n234_), .A2(KEYINPUT24), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n213_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n385_), .B1(new_n232_), .B2(new_n231_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n230_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n238_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n377_), .B1(new_n344_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n339_), .A2(new_n342_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n393_), .A2(new_n337_), .B1(new_n322_), .B2(new_n332_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n229_), .A2(new_n240_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n376_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n344_), .B2(new_n391_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n376_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n394_), .A2(new_n395_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n374_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n382_), .A2(new_n386_), .B1(new_n389_), .B2(new_n238_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n394_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n243_), .A2(new_n244_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n344_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n376_), .A2(new_n398_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n400_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(KEYINPUT95), .A3(new_n407_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT20), .B1(new_n394_), .B2(new_n410_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n412_), .A2(new_n344_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n376_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n407_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT95), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n409_), .A2(new_n418_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n408_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n423_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n374_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n373_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n311_), .A2(new_n430_), .A3(KEYINPUT96), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT96), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n262_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n373_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n362_), .A2(new_n369_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n352_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n370_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n306_), .A2(new_n426_), .A3(new_n439_), .A4(new_n429_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n300_), .B(new_n298_), .C1(KEYINPUT4), .C2(new_n297_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n266_), .B(new_n269_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n295_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n427_), .A2(new_n423_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n305_), .B2(KEYINPUT93), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n305_), .A2(KEYINPUT93), .A3(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n304_), .A2(new_n305_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n407_), .A2(KEYINPUT32), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n417_), .B2(new_n451_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n448_), .A2(new_n449_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n440_), .B1(new_n454_), .B2(new_n439_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n262_), .A2(new_n310_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n431_), .A2(new_n435_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G8gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT74), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G22gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n256_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G15gat), .A2(G22gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G1gat), .A2(G8gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n462_), .A2(new_n463_), .B1(KEYINPUT14), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n460_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n460_), .A2(new_n465_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n460_), .B(new_n465_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n468_), .A2(new_n471_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n471_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n474_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n480_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n472_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT75), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT76), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G141gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  AND3_X1   g290(.A1(new_n487_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n457_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G230gat), .ZN(new_n497_));
  INV_X1    g296(.A(G233gat), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT65), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT65), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(G106gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(KEYINPUT64), .ZN(new_n517_));
  OR2_X1    g316(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(KEYINPUT64), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G85gat), .ZN(new_n522_));
  INV_X1    g321(.A(G92gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(KEYINPUT9), .A3(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n525_), .A2(KEYINPUT9), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n515_), .A2(new_n521_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n511_), .A2(KEYINPUT66), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n508_), .A2(new_n510_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n246_), .A3(new_n516_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n524_), .A2(new_n525_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n530_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(KEYINPUT8), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n515_), .B2(new_n537_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n506_), .B(new_n529_), .C1(new_n541_), .C2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT67), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT65), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT65), .B1(new_n508_), .B2(new_n510_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n537_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n542_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n532_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n535_), .A2(new_n536_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n539_), .B1(new_n553_), .B2(new_n533_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n554_), .B2(new_n530_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n506_), .A4(new_n529_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n546_), .A2(KEYINPUT68), .A3(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n529_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n506_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT68), .B1(new_n546_), .B2(new_n557_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n499_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT12), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n547_), .A2(new_n548_), .ZN(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT64), .B(G106gat), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n518_), .A2(new_n519_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n527_), .B(new_n526_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT69), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n515_), .A2(new_n571_), .A3(new_n528_), .A4(new_n521_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n555_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n503_), .B(KEYINPUT12), .C1(new_n504_), .C2(new_n505_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n565_), .A2(new_n561_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n499_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n545_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G120gat), .B(G148gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G176gat), .B(G204gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n564_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n564_), .A2(new_n580_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n585_), .B(KEYINPUT71), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n586_), .B(new_n587_), .C1(new_n588_), .C2(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n564_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n564_), .B2(new_n580_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT13), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n506_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n474_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT17), .ZN(new_n600_));
  XOR2_X1   g399(.A(G127gat), .B(G155gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n599_), .A2(new_n600_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(KEYINPUT17), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n538_), .A2(new_n540_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n610_), .A2(KEYINPUT8), .B1(new_n549_), .B2(new_n542_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n570_), .A2(new_n572_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n473_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT35), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n555_), .A2(new_n471_), .A3(new_n529_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n616_), .A2(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n613_), .A2(new_n623_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT36), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT72), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n628_), .B(KEYINPUT36), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n625_), .B2(new_n634_), .ZN(new_n635_));
  AOI211_X1 g434(.A(KEYINPUT72), .B(new_n633_), .C1(new_n622_), .C2(new_n624_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n630_), .B(new_n631_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n625_), .A2(new_n629_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n633_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT37), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n609_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n596_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n496_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT97), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n496_), .A2(new_n646_), .A3(new_n643_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n265_), .A3(new_n450_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n635_), .A2(new_n636_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n630_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT98), .Z(new_n654_));
  INV_X1    g453(.A(new_n445_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n305_), .A2(KEYINPUT93), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT33), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n657_), .A3(new_n449_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n453_), .A2(new_n450_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n439_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AND4_X1   g459(.A1(new_n306_), .A2(new_n426_), .A3(new_n429_), .A4(new_n439_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n456_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT96), .B1(new_n311_), .B2(new_n430_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n433_), .A2(new_n434_), .A3(new_n432_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n662_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n654_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n596_), .A2(new_n495_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n608_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n265_), .B1(new_n668_), .B2(new_n450_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n651_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n650_), .B2(new_n649_), .ZN(G1324gat));
  NAND2_X1  g470(.A1(new_n426_), .A2(new_n429_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(G8gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n645_), .A2(new_n647_), .A3(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n666_), .A2(new_n667_), .A3(new_n672_), .A4(new_n608_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT39), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G8gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G8gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT100), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n675_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n681_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  INV_X1    g486(.A(new_n456_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n256_), .B1(new_n668_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n648_), .A2(new_n256_), .A3(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n439_), .A2(new_n461_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT103), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n648_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n668_), .A2(new_n439_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G22gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT102), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n699_), .A3(G22gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n701_));
  AND3_X1   g500(.A1(new_n698_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n695_), .B1(new_n702_), .B2(new_n703_), .ZN(G1327gat));
  NOR3_X1   g503(.A1(new_n596_), .A2(new_n495_), .A3(new_n608_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n637_), .A2(new_n640_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  INV_X1    g507(.A(new_n706_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n665_), .A2(KEYINPUT104), .A3(new_n708_), .A4(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n431_), .A2(new_n435_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n706_), .B1(new_n712_), .B2(new_n662_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT104), .B1(new_n713_), .B2(new_n708_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT44), .B(new_n705_), .C1(new_n711_), .C2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT105), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n665_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(new_n707_), .A3(new_n710_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(KEYINPUT44), .A4(new_n705_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n705_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n450_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G29gat), .B1(new_n724_), .B2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n652_), .A2(new_n609_), .A3(new_n630_), .ZN(new_n730_));
  NOR4_X1   g529(.A1(new_n457_), .A2(new_n495_), .A3(new_n596_), .A4(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n306_), .A2(G29gat), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT106), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n729_), .A2(new_n734_), .ZN(G1328gat));
  AOI21_X1  g534(.A(new_n673_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n723_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G36gat), .ZN(new_n738_));
  INV_X1    g537(.A(G36gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n731_), .A2(new_n739_), .A3(new_n672_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT45), .Z(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(KEYINPUT46), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n739_), .B1(new_n723_), .B2(new_n736_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n741_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1329gat));
  AND2_X1   g546(.A1(new_n731_), .A2(new_n688_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(G43gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n727_), .A2(G43gat), .A3(new_n688_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n724_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n749_), .B(new_n752_), .C1(new_n724_), .C2(new_n750_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1330gat));
  NAND2_X1  g555(.A1(new_n727_), .A2(new_n439_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G50gat), .B1(new_n724_), .B2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n373_), .A2(G50gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT108), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n731_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1331gat));
  NOR2_X1   g561(.A1(new_n595_), .A2(new_n494_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n457_), .A2(new_n642_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n450_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n654_), .ZN(new_n767_));
  NOR4_X1   g566(.A1(new_n767_), .A2(new_n457_), .A3(new_n609_), .A4(new_n764_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n306_), .A2(KEYINPUT109), .ZN(new_n769_));
  MUX2_X1   g568(.A(KEYINPUT109), .B(new_n769_), .S(G57gat), .Z(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n768_), .B2(new_n770_), .ZN(G1332gat));
  INV_X1    g570(.A(G64gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n768_), .B2(new_n672_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT48), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n765_), .A2(new_n772_), .A3(new_n672_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1333gat));
  INV_X1    g575(.A(G71gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n765_), .A2(new_n777_), .A3(new_n688_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n768_), .A2(new_n688_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G71gat), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT49), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT49), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n768_), .B2(new_n439_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT50), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n765_), .A2(new_n785_), .A3(new_n439_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n457_), .A2(new_n764_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n730_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT111), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n794_), .A3(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n522_), .A3(new_n450_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n764_), .A2(new_n608_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n720_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n450_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n801_), .B2(new_n522_), .ZN(G1336gat));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n523_), .A3(new_n672_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n672_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n805_), .B2(new_n523_), .ZN(G1337gat));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n456_), .A2(new_n568_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n796_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n796_), .B2(new_n808_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n720_), .A2(new_n688_), .A3(new_n798_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n246_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT113), .B(KEYINPUT51), .C1(new_n811_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n816_));
  OAI221_X1 g615(.A(new_n816_), .B1(new_n813_), .B2(new_n246_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1338gat));
  NOR2_X1   g617(.A1(new_n373_), .A2(new_n567_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n796_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT114), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n796_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n720_), .A2(new_n439_), .A3(new_n798_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(new_n516_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n824_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n824_), .A2(new_n828_), .A3(new_n832_), .A4(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n575_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n506_), .B1(new_n555_), .B2(new_n529_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(KEYINPUT12), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n838_), .B2(new_n578_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n561_), .A2(new_n565_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n579_), .A2(new_n840_), .A3(KEYINPUT55), .A4(new_n836_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n576_), .A2(new_n843_), .A3(new_n546_), .A4(new_n557_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n840_), .A2(new_n546_), .A3(new_n557_), .A4(new_n836_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n577_), .B1(new_n845_), .B2(KEYINPUT116), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n842_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n590_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n848_), .A2(new_n586_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n476_), .A2(new_n478_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n481_), .A2(new_n483_), .A3(new_n480_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  MUX2_X1   g651(.A(new_n852_), .B(new_n487_), .S(new_n491_), .Z(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n546_), .A2(new_n557_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT116), .B1(new_n838_), .B2(new_n855_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n844_), .A2(new_n499_), .A3(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n854_), .B(new_n589_), .C1(new_n857_), .C2(new_n842_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n849_), .A2(KEYINPUT58), .A3(new_n853_), .A4(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n848_), .A2(new_n586_), .A3(new_n853_), .A4(new_n858_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n706_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n859_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI211_X1 g663(.A(KEYINPUT118), .B(new_n706_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n848_), .A2(new_n494_), .A3(new_n586_), .A4(new_n858_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n853_), .B1(new_n593_), .B2(new_n592_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n653_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(KEYINPUT57), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n869_), .B(new_n653_), .C1(new_n871_), .C2(KEYINPUT57), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n609_), .B1(new_n866_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n595_), .A2(new_n641_), .A3(new_n877_), .A4(new_n495_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT115), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n595_), .A2(new_n641_), .A3(new_n495_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT54), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n878_), .A2(KEYINPUT115), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n876_), .A2(new_n885_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n434_), .A2(new_n456_), .A3(new_n306_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G113gat), .B1(new_n889_), .B2(new_n494_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n874_), .B(new_n873_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n609_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n609_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n885_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n887_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n888_), .A2(KEYINPUT59), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(G113gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n494_), .A2(KEYINPUT120), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(G113gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n890_), .B1(new_n902_), .B2(new_n906_), .ZN(G1340gat));
  OAI21_X1  g706(.A(G120gat), .B1(new_n901_), .B2(new_n595_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n595_), .A2(KEYINPUT60), .ZN(new_n909_));
  MUX2_X1   g708(.A(new_n909_), .B(KEYINPUT60), .S(G120gat), .Z(new_n910_));
  NAND2_X1  g709(.A1(new_n889_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(G1341gat));
  OAI21_X1  g711(.A(G127gat), .B1(new_n901_), .B2(new_n609_), .ZN(new_n913_));
  OR3_X1    g712(.A1(new_n888_), .A2(G127gat), .A3(new_n609_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1342gat));
  OAI21_X1  g714(.A(G134gat), .B1(new_n901_), .B2(new_n706_), .ZN(new_n916_));
  OR3_X1    g715(.A1(new_n888_), .A2(G134gat), .A3(new_n654_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1343gat));
  NOR4_X1   g717(.A1(new_n688_), .A2(new_n306_), .A3(new_n373_), .A4(new_n672_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n886_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n494_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n596_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g724(.A(KEYINPUT61), .B(G155gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT121), .B1(new_n920_), .B2(new_n609_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n920_), .A2(KEYINPUT121), .A3(new_n609_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n927_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n930_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(new_n928_), .A3(new_n926_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1346gat));
  AND3_X1   g733(.A1(new_n921_), .A2(G162gat), .A3(new_n709_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n920_), .A2(new_n654_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937_));
  OR3_X1    g736(.A1(new_n936_), .A2(new_n937_), .A3(G162gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n936_), .B2(G162gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n673_), .A2(new_n433_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n439_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n895_), .A2(new_n494_), .A3(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(G169gat), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n944_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n895_), .A2(new_n236_), .A3(new_n494_), .A4(new_n943_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(G1348gat));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n886_), .B2(new_n373_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n884_), .B1(new_n891_), .B2(new_n609_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n953_), .A2(KEYINPUT123), .A3(new_n439_), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n952_), .A2(new_n954_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n942_), .A2(new_n237_), .A3(new_n595_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n895_), .A2(new_n596_), .A3(new_n943_), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n955_), .A2(new_n956_), .B1(new_n237_), .B2(new_n957_), .ZN(G1349gat));
  NAND2_X1  g757(.A1(new_n379_), .A2(new_n381_), .ZN(new_n959_));
  AND4_X1   g758(.A1(new_n959_), .A2(new_n895_), .A3(new_n608_), .A4(new_n943_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n942_), .A2(new_n609_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n961_), .B1(new_n952_), .B2(new_n954_), .ZN(new_n962_));
  AOI21_X1  g761(.A(G183gat), .B1(new_n962_), .B2(KEYINPUT124), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n964_), .B(new_n961_), .C1(new_n952_), .C2(new_n954_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n960_), .B1(new_n963_), .B2(new_n965_), .ZN(G1350gat));
  NAND4_X1  g765(.A1(new_n895_), .A2(new_n216_), .A3(new_n767_), .A4(new_n943_), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n895_), .A2(new_n709_), .A3(new_n943_), .ZN(new_n968_));
  INV_X1    g767(.A(G190gat), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n967_), .B1(new_n968_), .B2(new_n969_), .ZN(G1351gat));
  XNOR2_X1  g769(.A(KEYINPUT126), .B(G197gat), .ZN(new_n971_));
  NOR4_X1   g770(.A1(new_n688_), .A2(new_n673_), .A3(new_n450_), .A4(new_n373_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n886_), .A2(new_n972_), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n886_), .A2(KEYINPUT125), .A3(new_n972_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n971_), .B1(new_n977_), .B2(new_n494_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n971_), .ZN(new_n979_));
  AOI211_X1 g778(.A(new_n495_), .B(new_n979_), .C1(new_n975_), .C2(new_n976_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n978_), .A2(new_n980_), .ZN(G1352gat));
  INV_X1    g780(.A(new_n976_), .ZN(new_n982_));
  AOI21_X1  g781(.A(KEYINPUT125), .B1(new_n886_), .B2(new_n972_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  OAI21_X1  g783(.A(G204gat), .B1(new_n984_), .B2(new_n595_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n977_), .A2(new_n312_), .A3(new_n596_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n985_), .A2(new_n986_), .ZN(G1353gat));
  OR2_X1    g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n988_), .B1(new_n977_), .B2(new_n608_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(KEYINPUT63), .B(G211gat), .ZN(new_n990_));
  AOI211_X1 g789(.A(new_n609_), .B(new_n990_), .C1(new_n975_), .C2(new_n976_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n989_), .A2(new_n991_), .ZN(G1354gat));
  OAI21_X1  g791(.A(G218gat), .B1(new_n984_), .B2(new_n706_), .ZN(new_n993_));
  NAND3_X1  g792(.A1(new_n977_), .A2(new_n326_), .A3(new_n767_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n993_), .A2(new_n994_), .ZN(G1355gat));
endmodule


