//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n204_));
  AND2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT1), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT88), .B1(new_n207_), .B2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n212_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n218_), .A2(new_n221_), .A3(new_n222_), .A4(new_n211_), .ZN(new_n223_));
  AND3_X1   g022(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT89), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT3), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(KEYINPUT89), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n205_), .A2(new_n206_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n214_), .A2(new_n223_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n204_), .B1(new_n233_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n214_), .A2(new_n223_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n232_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n234_), .B(new_n235_), .Z(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(new_n204_), .A3(new_n241_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n203_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n203_), .ZN(new_n256_));
  AOI211_X1 g055(.A(KEYINPUT96), .B(new_n202_), .C1(new_n252_), .C2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n203_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT96), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n255_), .A2(new_n251_), .A3(new_n203_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n245_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n249_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n258_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G190gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT82), .B(G183gat), .C1(new_n266_), .C2(KEYINPUT81), .ZN(new_n267_));
  NAND2_X1  g066(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT25), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT81), .B1(new_n266_), .B2(G183gat), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n265_), .A2(new_n267_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT24), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(G169gat), .B2(G176gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  INV_X1    g074(.A(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n272_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n272_), .A2(KEYINPUT84), .A3(new_n280_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(G183gat), .A3(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n278_), .A2(new_n279_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n273_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n283_), .A2(new_n284_), .A3(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G169gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n288_), .A2(KEYINPUT85), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(new_n286_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT91), .ZN(new_n301_));
  INV_X1    g100(.A(G218gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G211gat), .ZN(new_n303_));
  INV_X1    g102(.A(G211gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G218gat), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n303_), .A2(new_n305_), .A3(KEYINPUT90), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT90), .B1(new_n303_), .B2(new_n305_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G197gat), .A2(G204gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT21), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT21), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n301_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n304_), .A2(G218gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n302_), .A2(G211gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n303_), .A2(new_n305_), .A3(KEYINPUT90), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(KEYINPUT91), .A3(new_n312_), .A4(new_n315_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n314_), .A2(new_n309_), .A3(new_n313_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n326_), .A3(new_n322_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT92), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n321_), .A2(new_n326_), .A3(KEYINPUT92), .A4(new_n322_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n300_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT20), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n317_), .A2(new_n324_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n265_), .A2(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n291_), .A2(new_n337_), .A3(new_n280_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n287_), .B(new_n296_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n289_), .B1(G183gat), .B2(G190gat), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n338_), .A2(new_n339_), .B1(new_n340_), .B2(new_n295_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n334_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n338_), .A2(new_n339_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n340_), .A2(new_n295_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n334_), .B1(new_n332_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n345_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n335_), .A2(new_n299_), .A3(new_n293_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n346_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n300_), .A2(new_n332_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT20), .B1(new_n335_), .B2(new_n341_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n345_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n333_), .A2(new_n342_), .A3(new_n351_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT18), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n364_));
  MUX2_X1   g163(.A(new_n354_), .B(new_n359_), .S(new_n364_), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n264_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G22gat), .B(G50gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n233_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n233_), .B2(new_n370_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n368_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT28), .B1(new_n240_), .B2(KEYINPUT29), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT94), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n379_), .A3(new_n376_), .ZN(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n381_));
  OAI21_X1  g180(.A(new_n332_), .B1(new_n233_), .B2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(G228gat), .A2(G233gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n335_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n240_), .A2(KEYINPUT29), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n382_), .A2(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n378_), .A2(new_n380_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n382_), .A2(new_n383_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n384_), .A2(new_n385_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT94), .B(new_n377_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G78gat), .B(G106gat), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n392_), .A3(new_n390_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n258_), .A2(new_n398_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n245_), .A2(new_n398_), .A3(new_n249_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT97), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n203_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n202_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n404_), .A2(new_n263_), .A3(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n357_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n363_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT97), .B(new_n400_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n399_), .A2(new_n403_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n366_), .A2(new_n397_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT86), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT30), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G227gat), .A2(G233gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n417_), .B(G71gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G99gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n293_), .A2(new_n299_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n421_), .A2(new_n416_), .A3(new_n422_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n236_), .B(KEYINPUT31), .ZN(new_n426_));
  OR4_X1    g225(.A1(KEYINPUT87), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT87), .B1(new_n424_), .B2(new_n425_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n423_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n431_), .A3(new_n426_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n245_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n249_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n357_), .A2(new_n363_), .A3(new_n358_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT27), .B(new_n440_), .C1(new_n354_), .C2(new_n363_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n436_), .A2(new_n439_), .A3(new_n441_), .A4(new_n258_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n433_), .B1(new_n442_), .B2(new_n396_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n412_), .A2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n363_), .B1(new_n346_), .B2(new_n353_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n407_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n363_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n359_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n437_), .B1(new_n449_), .B2(new_n440_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT99), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n441_), .A2(new_n452_), .A3(new_n439_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n396_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n427_), .A2(new_n432_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n264_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n444_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT73), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G43gat), .B(G50gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n459_), .A2(KEYINPUT73), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(KEYINPUT73), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n463_), .A2(KEYINPUT15), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT15), .B1(new_n463_), .B2(new_n466_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT76), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT76), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n474_), .B(KEYINPUT14), .C1(new_n470_), .C2(new_n471_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n469_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n463_), .A2(new_n466_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n482_), .B(new_n479_), .Z(new_n486_));
  INV_X1    g285(.A(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT80), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n489_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT6), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT9), .ZN(new_n499_));
  OR2_X1    g298(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT9), .A3(new_n498_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n497_), .A2(new_n499_), .A3(new_n503_), .A4(new_n505_), .ZN(new_n506_));
  OR3_X1    g305(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n496_), .A2(KEYINPUT6), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n507_), .B(new_n508_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT8), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n504_), .A2(new_n498_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT66), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n513_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n506_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G71gat), .B(G78gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(KEYINPUT11), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n520_), .B2(KEYINPUT11), .ZN(new_n523_));
  INV_X1    g322(.A(G64gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G57gat), .ZN(new_n525_));
  INV_X1    g324(.A(G57gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G64gat), .ZN(new_n527_));
  AND4_X1   g326(.A1(new_n522_), .A2(new_n525_), .A3(new_n527_), .A4(KEYINPUT11), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n521_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n527_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT11), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT67), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n520_), .A2(new_n522_), .A3(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .A4(new_n519_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n518_), .A2(new_n536_), .A3(KEYINPUT12), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT12), .B1(new_n518_), .B2(new_n536_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n506_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n512_), .A2(new_n515_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT8), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n512_), .A2(new_n515_), .A3(new_n513_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n529_), .A2(new_n535_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n543_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n518_), .B2(new_n536_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(KEYINPUT68), .A3(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n518_), .A2(new_n536_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n539_), .A2(new_n550_), .B1(new_n555_), .B2(new_n543_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G120gat), .B(G148gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT71), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT69), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n561_), .B1(new_n556_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n555_), .A2(new_n543_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n538_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n518_), .A2(new_n536_), .A3(KEYINPUT12), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n550_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(KEYINPUT69), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n563_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n562_), .B1(new_n570_), .B2(KEYINPUT69), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n556_), .A2(new_n564_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(KEYINPUT71), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n572_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n495_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n570_), .B2(new_n561_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n565_), .A2(new_n571_), .A3(new_n580_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT13), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n572_), .A2(new_n576_), .A3(new_n575_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT72), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n494_), .B1(new_n579_), .B2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n458_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n479_), .B(new_n549_), .ZN(new_n589_));
  AND2_X1   g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n590_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n591_), .A2(KEYINPUT78), .A3(new_n593_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n603_), .A3(new_n601_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n468_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n463_), .A2(KEYINPUT15), .A3(new_n466_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n518_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT74), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n548_), .A2(new_n482_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n611_), .A2(new_n612_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT36), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n616_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n611_), .A2(new_n618_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n617_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n611_), .B2(KEYINPUT74), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n619_), .B(new_n623_), .C1(new_n626_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT75), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n629_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n612_), .B1(new_n469_), .B2(new_n518_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n625_), .B1(new_n635_), .B2(new_n627_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n636_), .B2(new_n619_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n631_), .B(KEYINPUT37), .C1(new_n632_), .C2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n619_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n633_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n640_), .B(new_n629_), .C1(new_n630_), .C2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n608_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT79), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n588_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n470_), .A3(new_n264_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n587_), .A2(new_n608_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n412_), .A2(new_n443_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n632_), .A2(new_n637_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n264_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G1gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n648_), .A2(new_n649_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n650_), .A2(new_n656_), .A3(new_n657_), .ZN(G1324gat));
  NAND2_X1  g457(.A1(new_n451_), .A2(new_n453_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n651_), .A2(new_n660_), .A3(new_n654_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(KEYINPUT100), .A3(G8gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT100), .B1(new_n661_), .B2(G8gat), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n647_), .A2(new_n471_), .A3(new_n660_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT40), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1325gat));
  NAND3_X1  g472(.A1(new_n651_), .A2(new_n433_), .A3(new_n654_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G15gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT101), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT41), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT41), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n646_), .A2(G15gat), .A3(new_n455_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT102), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n678_), .A3(new_n680_), .ZN(G1326gat));
  NAND3_X1  g480(.A1(new_n651_), .A2(new_n396_), .A3(new_n654_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(G22gat), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G22gat), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n397_), .A2(G22gat), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n684_), .A2(new_n685_), .B1(new_n646_), .B2(new_n686_), .ZN(G1327gat));
  NAND2_X1  g486(.A1(new_n607_), .A2(new_n653_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n588_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n264_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n587_), .A2(new_n607_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n638_), .A2(new_n642_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n458_), .B2(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n652_), .A2(KEYINPUT43), .A3(new_n643_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n693_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n264_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n692_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n660_), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G36gat), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT105), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n659_), .A2(G36gat), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n458_), .A2(new_n690_), .A3(new_n587_), .A4(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n711_), .A2(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(KEYINPUT45), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n712_), .A2(new_n713_), .B1(KEYINPUT105), .B2(new_n707_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n706_), .A2(new_n709_), .A3(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n709_), .B1(new_n706_), .B2(new_n714_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  AND2_X1   g516(.A1(new_n433_), .A2(G43gat), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n700_), .A2(new_n701_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G43gat), .B1(new_n691_), .B2(new_n433_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n691_), .B2(new_n396_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n396_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n702_), .B2(new_n727_), .ZN(G1331gat));
  NAND2_X1  g527(.A1(new_n579_), .A2(new_n586_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n494_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n645_), .A2(new_n458_), .A3(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n526_), .A3(new_n264_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n729_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n605_), .A2(new_n606_), .A3(new_n494_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n654_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n264_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G57gat), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n733_), .A2(new_n739_), .ZN(G1332gat));
  NAND3_X1  g539(.A1(new_n732_), .A2(new_n524_), .A3(new_n660_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  INV_X1    g541(.A(new_n737_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n660_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(G64gat), .ZN(new_n745_));
  AOI211_X1 g544(.A(KEYINPUT48), .B(new_n524_), .C1(new_n743_), .C2(new_n660_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n745_), .B2(new_n746_), .ZN(G1333gat));
  NOR2_X1   g546(.A1(new_n455_), .A2(G71gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT107), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n732_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G71gat), .B1(new_n737_), .B2(new_n455_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT49), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT49), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1334gat));
  INV_X1    g553(.A(G78gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n732_), .A2(new_n755_), .A3(new_n396_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n743_), .A2(new_n396_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(G78gat), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G78gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1335gat));
  AND3_X1   g560(.A1(new_n731_), .A2(new_n458_), .A3(new_n690_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n264_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n696_), .A2(new_n697_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n730_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n579_), .A2(new_n586_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n579_), .A2(new_n586_), .A3(KEYINPUT109), .A4(new_n765_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n264_), .A2(G85gat), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT110), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n770_), .B2(new_n772_), .ZN(G1336gat));
  INV_X1    g572(.A(G92gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n762_), .A2(new_n774_), .A3(new_n660_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n770_), .A2(new_n660_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n774_), .ZN(G1337gat));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n778_), .A2(KEYINPUT51), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n768_), .A2(new_n769_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n433_), .B(new_n780_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G99gat), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n433_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n762_), .A2(KEYINPUT112), .A3(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n731_), .A2(new_n690_), .A3(new_n458_), .A4(new_n785_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n786_), .A2(new_n789_), .B1(new_n778_), .B2(KEYINPUT51), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n779_), .B1(new_n784_), .B2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n782_), .A2(new_n783_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT111), .B1(new_n781_), .B2(G99gat), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n779_), .B(new_n790_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n791_), .A2(new_n795_), .ZN(G1338gat));
  OAI211_X1 g595(.A(new_n396_), .B(new_n780_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G106gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT115), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(new_n800_), .A3(G106gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(KEYINPUT52), .A3(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n397_), .A2(G106gat), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n731_), .A2(new_n690_), .A3(new_n458_), .A4(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT114), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n800_), .B1(new_n797_), .B2(G106gat), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n802_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n802_), .B2(new_n808_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1339gat));
  NOR2_X1   g611(.A1(new_n695_), .A2(new_n735_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n577_), .A2(new_n578_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n815_), .B2(KEYINPUT54), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n813_), .A2(new_n818_), .A3(new_n814_), .A4(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n816_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT122), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n493_), .B1(new_n486_), .B2(new_n484_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n480_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n485_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n570_), .A2(new_n561_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n539_), .A2(KEYINPUT55), .A3(new_n550_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n569_), .A2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n539_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n830_), .B(new_n832_), .C1(new_n833_), .C2(new_n542_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n561_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n829_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n643_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n836_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(KEYINPUT58), .A4(new_n829_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT58), .B(new_n829_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT119), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n839_), .A2(new_n844_), .A3(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n494_), .A2(new_n828_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n836_), .B2(new_n835_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n572_), .A2(new_n575_), .A3(new_n826_), .A4(new_n825_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n653_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n822_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(KEYINPUT57), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n839_), .A2(new_n844_), .A3(new_n846_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(KEYINPUT122), .C1(new_n851_), .C2(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n821_), .B1(new_n858_), .B2(new_n607_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n738_), .A2(new_n455_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n454_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT120), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n856_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n855_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n607_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n816_), .A2(new_n817_), .A3(new_n820_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n862_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n859_), .A2(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G113gat), .B1(new_n871_), .B2(new_n494_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n869_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n494_), .A2(G113gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(G120gat), .B1(new_n871_), .B2(new_n729_), .ZN(new_n876_));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(KEYINPUT60), .B2(new_n877_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n876_), .B1(new_n873_), .B2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n871_), .B2(new_n607_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n607_), .A2(G127gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n873_), .B2(new_n882_), .ZN(G1342gat));
  OAI21_X1  g682(.A(G134gat), .B1(new_n871_), .B2(new_n643_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n632_), .A2(new_n637_), .A3(G134gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n873_), .B2(new_n885_), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n867_), .A2(new_n868_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n397_), .A2(new_n433_), .ZN(new_n888_));
  AND4_X1   g687(.A1(new_n659_), .A2(new_n887_), .A3(new_n264_), .A4(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n730_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n734_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n608_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n889_), .A2(new_n897_), .A3(new_n653_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n889_), .A2(new_n695_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1347gat));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n660_), .A2(new_n397_), .A3(new_n456_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n859_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n866_), .B1(new_n865_), .B2(new_n822_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n608_), .B1(new_n905_), .B2(new_n857_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT123), .B(new_n904_), .C1(new_n906_), .C2(new_n821_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT22), .B(G169gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n730_), .A2(new_n909_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT124), .Z(new_n911_));
  NAND2_X1  g710(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n730_), .B(new_n904_), .C1(new_n906_), .C2(new_n821_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n913_), .A2(new_n914_), .A3(G169gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n913_), .B2(G169gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n912_), .B1(new_n915_), .B2(new_n916_), .ZN(G1348gat));
  INV_X1    g716(.A(new_n887_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n918_), .A2(new_n277_), .A3(new_n729_), .A4(new_n902_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n908_), .A2(new_n734_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n277_), .ZN(G1349gat));
  NOR2_X1   g720(.A1(new_n918_), .A2(new_n902_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G183gat), .B1(new_n922_), .B2(new_n608_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n607_), .A2(new_n336_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n908_), .B2(new_n924_), .ZN(G1350gat));
  AND2_X1   g724(.A1(new_n653_), .A2(new_n265_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n908_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(G190gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n643_), .B1(new_n903_), .B2(new_n907_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1351gat));
  NAND2_X1  g729(.A1(new_n888_), .A2(new_n738_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT125), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n932_), .A2(new_n660_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n887_), .A2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n887_), .A2(KEYINPUT126), .A3(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938_), .B2(new_n730_), .ZN(new_n939_));
  INV_X1    g738(.A(G197gat), .ZN(new_n940_));
  AOI211_X1 g739(.A(new_n940_), .B(new_n494_), .C1(new_n936_), .C2(new_n937_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1352gat));
  INV_X1    g741(.A(new_n937_), .ZN(new_n943_));
  AOI21_X1  g742(.A(KEYINPUT126), .B1(new_n887_), .B2(new_n933_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n734_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n945_), .A2(KEYINPUT127), .A3(G204gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n938_), .A2(new_n734_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1353gat));
  OR2_X1    g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n950_), .B1(new_n938_), .B2(new_n608_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT63), .B(G211gat), .ZN(new_n952_));
  AOI211_X1 g751(.A(new_n607_), .B(new_n952_), .C1(new_n936_), .C2(new_n937_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1354gat));
  NAND3_X1  g753(.A1(new_n938_), .A2(new_n302_), .A3(new_n653_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n643_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n302_), .B2(new_n956_), .ZN(G1355gat));
endmodule


