//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  AND2_X1   g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n204_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n203_), .A3(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G183gat), .ZN(new_n226_));
  INV_X1    g025(.A(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n209_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n221_), .A2(new_n218_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n216_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n232_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n238_), .A3(KEYINPUT82), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n215_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G99gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(G43gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n243_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n249_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G227gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(G15gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT30), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT31), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n257_), .A3(new_n251_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n262_));
  INV_X1    g061(.A(G155gat), .ZN(new_n263_));
  INV_X1    g062(.A(G162gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT85), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(KEYINPUT85), .A3(G155gat), .A4(G162gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n267_), .A2(new_n269_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G141gat), .ZN(new_n275_));
  INV_X1    g074(.A(G148gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT83), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(G141gat), .B2(G148gat), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n277_), .A2(new_n279_), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n282_), .A2(new_n285_), .A3(new_n286_), .A4(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n265_), .A2(new_n266_), .B1(G155gat), .B2(G162gat), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n274_), .A2(new_n280_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT29), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G22gat), .B(G50gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT28), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n292_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G78gat), .B(G106gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G228gat), .A2(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n274_), .A2(new_n280_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n289_), .A2(new_n288_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n291_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G197gat), .A2(G204gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G197gat), .A2(G204gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(KEYINPUT21), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n308_), .A2(new_n309_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n299_), .B1(new_n302_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n311_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n298_), .B(new_n314_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n297_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n295_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n278_), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT83), .B1(new_n275_), .B2(new_n276_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n283_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n265_), .A2(new_n266_), .B1(KEYINPUT1), .B2(new_n268_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n271_), .A2(new_n273_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n301_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT29), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n298_), .B1(new_n326_), .B2(new_n314_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n315_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n296_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n313_), .A2(new_n315_), .A3(new_n297_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n318_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n329_), .A2(new_n295_), .A3(new_n317_), .A4(new_n330_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G85gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT0), .B(G57gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n290_), .B2(new_n249_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n247_), .A2(new_n248_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n247_), .A2(new_n248_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n341_), .B(new_n344_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT87), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n300_), .A2(new_n301_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(new_n341_), .A3(new_n339_), .A4(new_n344_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n344_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n290_), .A2(new_n249_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n347_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n338_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n354_), .A3(new_n338_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n261_), .A2(new_n334_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT97), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n234_), .B1(new_n361_), .B2(new_n209_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT24), .B1(new_n221_), .B2(new_n218_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n240_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n222_), .A2(new_n231_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n242_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n212_), .A2(new_n214_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n204_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n312_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n216_), .A2(new_n203_), .A3(new_n220_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n208_), .A2(new_n211_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n213_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n373_));
  OAI22_X1  g172(.A1(new_n232_), .A2(new_n372_), .B1(new_n373_), .B2(new_n204_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n314_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n370_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n366_), .A2(new_n369_), .A3(new_n312_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n374_), .B2(new_n314_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n379_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G8gat), .B(G36gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n378_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n372_), .ZN(new_n392_));
  OR2_X1    g191(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n393_));
  NAND2_X1  g192(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n205_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n214_), .B1(new_n395_), .B2(new_n234_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n365_), .A2(new_n392_), .B1(new_n396_), .B2(new_n368_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n381_), .B1(new_n397_), .B2(new_n312_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n243_), .B2(new_n312_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n377_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n380_), .A2(new_n382_), .A3(new_n379_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT93), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n380_), .A2(new_n382_), .A3(new_n403_), .A4(new_n379_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n387_), .B(KEYINPUT94), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n388_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n380_), .A2(new_n382_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n377_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n398_), .B(new_n379_), .C1(new_n243_), .C2(new_n312_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n387_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n391_), .A2(new_n408_), .B1(new_n414_), .B2(new_n390_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n359_), .A2(new_n360_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n360_), .B1(new_n359_), .B2(new_n415_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n387_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n390_), .B1(new_n389_), .B2(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n399_), .A2(new_n377_), .B1(new_n401_), .B2(KEYINPUT93), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n421_), .B2(new_n404_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n413_), .A2(KEYINPUT27), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n357_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(new_n355_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n334_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT95), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n358_), .B1(new_n333_), .B2(new_n332_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT95), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n415_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n334_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n389_), .A2(new_n419_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n346_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT91), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n346_), .A2(KEYINPUT91), .A3(new_n347_), .A4(new_n350_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n352_), .A2(new_n353_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n338_), .B1(new_n440_), .B2(new_n348_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT90), .B(KEYINPUT33), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n357_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n434_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n351_), .A2(KEYINPUT33), .A3(new_n354_), .A4(new_n338_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT92), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n444_), .A2(new_n413_), .A3(new_n409_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n446_), .B(KEYINPUT89), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .A4(new_n442_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n405_), .A2(KEYINPUT32), .A3(new_n387_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n378_), .A2(new_n383_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT32), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n388_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n358_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n432_), .B1(new_n433_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n261_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT96), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n433_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n428_), .A2(new_n431_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT96), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n261_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n418_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G229gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT74), .B(G8gat), .ZN(new_n470_));
  INV_X1    g269(.A(G1gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT75), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G8gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G43gat), .B(G50gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n476_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n475_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n469_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT77), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n480_), .B(KEYINPUT15), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n489_), .A3(new_n469_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G113gat), .B(G141gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G169gat), .B(G197gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT78), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(new_n497_), .A3(new_n490_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT79), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(KEYINPUT79), .A3(new_n498_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT98), .B1(new_n468_), .B2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n416_), .A2(new_n417_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n466_), .B1(new_n465_), .B2(new_n261_), .ZN(new_n506_));
  AOI211_X1 g305(.A(KEYINPUT96), .B(new_n461_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(new_n502_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT67), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT7), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT67), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G85gat), .B(G92gat), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT68), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(new_n529_), .A3(new_n526_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(KEYINPUT8), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n519_), .B(KEYINPUT66), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n522_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n526_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT10), .B(G99gat), .Z(new_n537_));
  INV_X1    g336(.A(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT64), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT64), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n537_), .A2(new_n541_), .A3(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n526_), .A2(KEYINPUT9), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT65), .B(G92gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(G85gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n532_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n536_), .B1(new_n544_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT69), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n552_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT66), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n519_), .B(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(new_n549_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n531_), .A2(new_n535_), .B1(new_n543_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(G230gat), .A2(G233gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n531_), .A2(new_n535_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n551_), .B2(new_n544_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(KEYINPUT70), .A3(new_n543_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(KEYINPUT12), .B(new_n561_), .C1(new_n571_), .C2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT12), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n566_), .B2(new_n560_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n569_), .B1(new_n566_), .B2(new_n560_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n570_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n570_), .A2(new_n580_), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(KEYINPUT71), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n581_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(KEYINPUT13), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT13), .B1(new_n589_), .B2(new_n591_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n514_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n591_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(KEYINPUT72), .A3(new_n592_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(KEYINPUT73), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(KEYINPUT73), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n560_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n483_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT17), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n611_), .B(KEYINPUT17), .Z(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n606_), .B2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n488_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT34), .ZN(new_n618_));
  OAI221_X1 g417(.A(new_n616_), .B1(KEYINPUT35), .B2(new_n618_), .C1(new_n484_), .C2(new_n552_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n619_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT36), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n619_), .B(new_n622_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n627_), .B(KEYINPUT36), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(KEYINPUT37), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n615_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n513_), .A2(new_n603_), .A3(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n471_), .A3(new_n358_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n639_), .A2(new_n644_), .A3(new_n640_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n600_), .A2(new_n499_), .A3(new_n615_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n633_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n468_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n600_), .A2(KEYINPUT100), .A3(new_n499_), .A4(new_n615_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n426_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n643_), .A2(new_n647_), .A3(new_n655_), .ZN(G1324gat));
  NAND3_X1  g455(.A1(new_n638_), .A2(new_n424_), .A3(new_n470_), .ZN(new_n657_));
  INV_X1    g456(.A(G8gat), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n654_), .A2(new_n415_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(KEYINPUT102), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n654_), .B2(new_n415_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n657_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n657_), .B(new_n667_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n654_), .B2(new_n261_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT105), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n674_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n638_), .A2(new_n254_), .A3(new_n461_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n654_), .B2(new_n433_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT42), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n433_), .A2(G22gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT106), .Z(new_n682_));
  NAND2_X1  g481(.A1(new_n638_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n633_), .A2(new_n615_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n600_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n504_), .B2(new_n511_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n358_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n634_), .A2(new_n636_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n468_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n634_), .A2(new_n636_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n508_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n615_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n600_), .A2(new_n499_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AND4_X1   g496(.A1(KEYINPUT107), .A2(new_n694_), .A3(KEYINPUT44), .A4(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT107), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(KEYINPUT44), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n358_), .A2(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n688_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n415_), .A2(G36gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n687_), .A2(KEYINPUT108), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT108), .B1(new_n687_), .B2(new_n709_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n686_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n512_), .A2(new_n714_), .A3(new_n709_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT45), .A3(new_n710_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n718_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n468_), .A2(KEYINPUT43), .A3(new_n689_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n691_), .B1(new_n508_), .B2(new_n692_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n697_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n415_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n706_), .B(new_n707_), .C1(new_n719_), .C2(new_n726_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n717_), .A2(KEYINPUT45), .A3(new_n710_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT45), .B1(new_n717_), .B2(new_n710_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n424_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n694_), .A2(KEYINPUT44), .A3(new_n697_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n699_), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G36gat), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n728_), .A2(new_n729_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT46), .B1(new_n737_), .B2(KEYINPUT109), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n727_), .A2(new_n738_), .ZN(G1329gat));
  NAND2_X1  g538(.A1(new_n461_), .A2(G43gat), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n701_), .A2(new_n702_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G43gat), .B1(new_n687_), .B2(new_n461_), .ZN(new_n742_));
  OR3_X1    g541(.A1(new_n741_), .A2(KEYINPUT47), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT47), .B1(new_n741_), .B2(new_n742_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1330gat));
  NOR3_X1   g544(.A1(new_n701_), .A2(new_n433_), .A3(new_n702_), .ZN(new_n746_));
  INV_X1    g545(.A(G50gat), .ZN(new_n747_));
  INV_X1    g546(.A(new_n687_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n334_), .A2(new_n747_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT110), .Z(new_n750_));
  OAI22_X1  g549(.A1(new_n746_), .A2(new_n747_), .B1(new_n748_), .B2(new_n750_), .ZN(G1331gat));
  NOR2_X1   g550(.A1(new_n600_), .A2(new_n637_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT111), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n468_), .A2(new_n499_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n358_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(KEYINPUT112), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT112), .B1(new_n755_), .B2(new_n756_), .ZN(new_n759_));
  NOR4_X1   g558(.A1(new_n601_), .A2(new_n602_), .A3(new_n510_), .A4(new_n695_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n652_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT113), .B(G57gat), .Z(new_n762_));
  NAND2_X1  g561(.A1(new_n358_), .A2(new_n762_), .ZN(new_n763_));
  OAI22_X1  g562(.A1(new_n758_), .A2(new_n759_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT114), .ZN(G1332gat));
  OAI21_X1  g564(.A(G64gat), .B1(new_n761_), .B2(new_n415_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT48), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n753_), .A2(new_n754_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n415_), .A2(G64gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT115), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n768_), .B2(new_n770_), .ZN(G1333gat));
  OAI21_X1  g570(.A(G71gat), .B1(new_n761_), .B2(new_n261_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT49), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n261_), .A2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n768_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n761_), .B2(new_n433_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT50), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n433_), .A2(G78gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n768_), .B2(new_n778_), .ZN(G1335gat));
  NOR4_X1   g578(.A1(new_n601_), .A2(new_n602_), .A3(new_n633_), .A4(new_n615_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n754_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(G85gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n358_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n694_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n600_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n499_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n695_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n785_), .A2(new_n426_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n784_), .B1(new_n783_), .B2(new_n789_), .ZN(G1336gat));
  AOI21_X1  g589(.A(G92gat), .B1(new_n782_), .B2(new_n424_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n785_), .A2(new_n788_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n424_), .A2(new_n546_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(G1337gat));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n461_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n795_), .A2(KEYINPUT116), .A3(G99gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT116), .B1(new_n795_), .B2(G99gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n461_), .A2(new_n537_), .ZN(new_n798_));
  OAI22_X1  g597(.A1(new_n796_), .A2(new_n797_), .B1(new_n781_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801_));
  OAI221_X1 g600(.A(new_n801_), .B1(new_n781_), .B2(new_n798_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1338gat));
  AOI21_X1  g602(.A(new_n538_), .B1(new_n792_), .B2(new_n334_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n780_), .A2(new_n538_), .A3(new_n334_), .A4(new_n754_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n805_), .A2(new_n808_), .A3(new_n812_), .A4(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n637_), .A2(new_n510_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n593_), .A2(new_n594_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NOR4_X1   g618(.A1(new_n637_), .A2(new_n510_), .A3(KEYINPUT54), .A4(new_n817_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n588_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n491_), .A2(new_n494_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n494_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n469_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n481_), .A2(new_n489_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n823_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n558_), .A2(new_n559_), .A3(KEYINPUT12), .ZN(new_n830_));
  INV_X1    g629(.A(new_n574_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT70), .B1(new_n565_), .B2(new_n543_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(new_n536_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n562_), .B2(new_n577_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n579_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n580_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n576_), .A2(new_n578_), .A3(new_n567_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n838_), .A2(new_n580_), .B1(new_n841_), .B2(new_n569_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n840_), .A2(KEYINPUT119), .A3(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n585_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n840_), .A2(KEYINPUT119), .A3(new_n842_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT119), .B1(new_n840_), .B2(new_n842_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT56), .B(new_n585_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n829_), .B1(new_n848_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n689_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(KEYINPUT58), .B(new_n829_), .C1(new_n848_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n498_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n497_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n588_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n585_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n863_), .B2(new_n851_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n596_), .B1(new_n828_), .B2(new_n823_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n633_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT57), .B(new_n633_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n857_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n821_), .B1(new_n870_), .B2(new_n695_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n415_), .A2(new_n358_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n261_), .A3(new_n334_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G113gat), .B1(new_n875_), .B2(new_n499_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(KEYINPUT120), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n855_), .A2(new_n856_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n615_), .B1(new_n883_), .B2(new_n869_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n873_), .B(new_n882_), .C1(new_n884_), .C2(new_n821_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n878_), .A2(new_n879_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n879_), .B1(new_n878_), .B2(new_n885_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n510_), .A2(G113gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n876_), .B1(new_n888_), .B2(new_n889_), .ZN(G1340gat));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n600_), .B2(KEYINPUT60), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n875_), .B(new_n892_), .C1(KEYINPUT60), .C2(new_n891_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n878_), .A2(new_n603_), .A3(new_n885_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n891_), .ZN(G1341gat));
  AOI21_X1  g694(.A(G127gat), .B1(new_n875_), .B2(new_n615_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n615_), .A2(G127gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n888_), .B2(new_n897_), .ZN(G1342gat));
  AOI21_X1  g697(.A(G134gat), .B1(new_n875_), .B2(new_n651_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n692_), .A2(G134gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n888_), .B2(new_n900_), .ZN(G1343gat));
  NOR2_X1   g700(.A1(new_n871_), .A2(new_n461_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n902_), .A2(new_n334_), .A3(new_n358_), .A4(new_n415_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT122), .B(G141gat), .Z(new_n904_));
  OR3_X1    g703(.A1(new_n903_), .A2(new_n787_), .A3(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n903_), .B2(new_n787_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1344gat));
  INV_X1    g706(.A(new_n603_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n903_), .A2(G148gat), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G148gat), .B1(new_n903_), .B2(new_n908_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1345gat));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n903_), .A2(new_n695_), .A3(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n695_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n903_), .B2(new_n689_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n651_), .A2(new_n264_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n903_), .B2(new_n917_), .ZN(G1347gat));
  NAND2_X1  g717(.A1(new_n359_), .A2(new_n424_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n499_), .B(new_n920_), .C1(new_n884_), .C2(new_n821_), .ZN(new_n921_));
  AOI21_X1  g720(.A(KEYINPUT123), .B1(new_n921_), .B2(G169gat), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n921_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(KEYINPUT62), .A3(new_n924_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT22), .B(G169gat), .Z(new_n926_));
  NOR2_X1   g725(.A1(new_n921_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n922_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n929_), .ZN(G1348gat));
  NOR2_X1   g729(.A1(new_n871_), .A2(new_n919_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G176gat), .B1(new_n932_), .B2(new_n908_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n220_), .A3(new_n786_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1349gat));
  OAI211_X1 g734(.A(new_n224_), .B(new_n226_), .C1(KEYINPUT124), .C2(G183gat), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n931_), .A2(new_n615_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n223_), .A2(KEYINPUT124), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n931_), .B2(new_n615_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n938_), .B2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n940_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n942_), .A2(new_n943_), .A3(new_n937_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n941_), .A2(new_n944_), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n932_), .B2(new_n689_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n651_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT126), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n932_), .B2(new_n948_), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n415_), .A2(new_n427_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n902_), .A2(new_n499_), .A3(new_n950_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g751(.A1(new_n902_), .A2(new_n603_), .A3(new_n950_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(KEYINPUT127), .B(G204gat), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1353gat));
  XNOR2_X1  g754(.A(KEYINPUT63), .B(G211gat), .ZN(new_n956_));
  OR2_X1    g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n902_), .A2(new_n615_), .A3(new_n950_), .ZN(new_n958_));
  MUX2_X1   g757(.A(new_n956_), .B(new_n957_), .S(new_n958_), .Z(G1354gat));
  NAND2_X1  g758(.A1(new_n902_), .A2(new_n950_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G218gat), .B1(new_n960_), .B2(new_n689_), .ZN(new_n961_));
  OR2_X1    g760(.A1(new_n633_), .A2(G218gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n960_), .B2(new_n962_), .ZN(G1355gat));
endmodule


