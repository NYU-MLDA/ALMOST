//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  INV_X1    g000(.A(G134gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G127gat), .ZN(new_n203_));
  INV_X1    g002(.A(G127gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G113gat), .ZN(new_n208_));
  INV_X1    g007(.A(G113gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G120gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT85), .B1(new_n206_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n211_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n203_), .A2(new_n205_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n212_), .B1(new_n215_), .B2(KEYINPUT85), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT31), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT86), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(G169gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT83), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n222_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n232_), .A2(new_n233_), .A3(G183gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n221_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n228_), .A2(KEYINPUT23), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n237_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT24), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n232_), .A2(new_n233_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(G190gat), .ZN(new_n251_));
  INV_X1    g050(.A(G183gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT25), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G183gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n248_), .B1(new_n250_), .B2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT26), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT25), .B(G183gat), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(KEYINPUT80), .A3(new_n261_), .A4(new_n251_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n247_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n244_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  AOI211_X1 g064(.A(KEYINPUT82), .B(new_n247_), .C1(new_n257_), .C2(new_n262_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n235_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G227gat), .A2(G233gat), .ZN(new_n268_));
  INV_X1    g067(.A(G15gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272_));
  INV_X1    g071(.A(G43gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n270_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n235_), .B(new_n276_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n271_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n275_), .B1(new_n271_), .B2(new_n277_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n219_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n219_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n278_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n218_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  NOR3_X1   g093(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n293_), .B(new_n294_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT3), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n290_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n303_));
  AND2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n298_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(KEYINPUT1), .B2(new_n289_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n215_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT98), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n216_), .A2(new_n307_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT98), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n302_), .A2(new_n311_), .A3(new_n306_), .A4(new_n215_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n309_), .A2(KEYINPUT4), .A3(new_n310_), .A4(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT4), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n216_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G225gat), .A2(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .A4(new_n316_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G1gat), .B(G29gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n321_), .A2(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n313_), .A2(new_n318_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT102), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n326_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT102), .B1(new_n333_), .B2(new_n319_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n328_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n217_), .A2(KEYINPUT86), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n281_), .A2(new_n284_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n286_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT94), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n239_), .A2(new_n238_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n230_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n222_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n344_), .B(new_n342_), .C1(new_n345_), .C2(new_n228_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT94), .ZN(new_n347_));
  INV_X1    g146(.A(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT26), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n261_), .A2(new_n251_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n246_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n245_), .A2(KEYINPUT93), .A3(KEYINPUT24), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n352_), .A2(new_n242_), .A3(new_n241_), .A4(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n343_), .A2(new_n347_), .A3(new_n350_), .A4(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G197gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(G204gat), .ZN(new_n357_));
  INV_X1    g156(.A(G204gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n358_), .A2(G197gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT21), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G211gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(G218gat), .ZN(new_n362_));
  INV_X1    g161(.A(G218gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(G211gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n356_), .B2(G204gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n356_), .A2(G204gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n358_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n360_), .B(new_n365_), .C1(new_n370_), .C2(KEYINPUT21), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT90), .B1(new_n362_), .B2(new_n364_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n363_), .A2(G211gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n361_), .A2(G218gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT90), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n372_), .A2(new_n370_), .A3(KEYINPUT21), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n221_), .B1(new_n237_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n355_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n382_), .A2(KEYINPUT20), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT96), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(KEYINPUT91), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n371_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n267_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n388_), .B1(new_n267_), .B2(new_n393_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n387_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n354_), .B(new_n350_), .C1(new_n346_), .C2(KEYINPUT94), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n341_), .B1(new_n230_), .B2(new_n342_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n381_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n378_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n403_), .B1(new_n407_), .B2(KEYINPUT95), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n392_), .B(new_n235_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n410_), .A3(new_n378_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n385_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n396_), .A2(new_n402_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n402_), .B1(new_n396_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n340_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n396_), .A2(new_n402_), .A3(new_n413_), .ZN(new_n417_));
  AND4_X1   g216(.A1(new_n386_), .A2(new_n408_), .A3(new_n409_), .A4(new_n411_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n382_), .A2(KEYINPUT20), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n420_), .B2(new_n385_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT27), .B(new_n417_), .C1(new_n421_), .C2(new_n402_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n307_), .A2(KEYINPUT29), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n378_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(G228gat), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G78gat), .B(G106gat), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n423_), .A2(new_n389_), .A3(new_n391_), .A4(new_n428_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT28), .B1(new_n307_), .B2(KEYINPUT29), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT28), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n302_), .A2(new_n438_), .A3(new_n439_), .A4(new_n306_), .ZN(new_n440_));
  XOR2_X1   g239(.A(G22gat), .B(G50gat), .Z(new_n441_));
  AND3_X1   g240(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n441_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n443_));
  OAI22_X1  g242(.A1(new_n435_), .A2(new_n436_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n436_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n443_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n434_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n416_), .A2(new_n422_), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n339_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n448_), .A2(new_n335_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n416_), .A2(new_n422_), .A3(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n412_), .A2(new_n385_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n387_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n267_), .A2(new_n393_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT96), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n267_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n401_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT100), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT100), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(new_n460_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n329_), .A2(new_n331_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .A4(new_n317_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n327_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n313_), .A2(new_n316_), .A3(new_n315_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT101), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n313_), .A2(KEYINPUT101), .A3(new_n316_), .A4(new_n315_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(KEYINPUT33), .A2(new_n466_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n459_), .A2(new_n465_), .A3(new_n417_), .A4(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n396_), .A2(new_n475_), .A3(new_n413_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n335_), .B(new_n476_), .C1(new_n421_), .C2(new_n475_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n448_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n452_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n286_), .A2(new_n338_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n450_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT75), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n486_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT76), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n490_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G36gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G29gat), .ZN(new_n495_));
  INV_X1    g294(.A(G29gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G36gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n273_), .A2(G50gat), .ZN(new_n498_));
  INV_X1    g297(.A(G50gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(G43gat), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n495_), .B(new_n497_), .C1(new_n498_), .C2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n497_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n493_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n493_), .A2(new_n508_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n501_), .A2(new_n504_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n505_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(KEYINPUT15), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n493_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n510_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G169gat), .B(G197gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n512_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n482_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT6), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G99gat), .A3(G106gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT10), .B(G99gat), .Z(new_n538_));
  INV_X1    g337(.A(G106gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT9), .ZN(new_n542_));
  INV_X1    g341(.A(G85gat), .ZN(new_n543_));
  INV_X1    g342(.A(G92gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT9), .A3(new_n541_), .ZN(new_n546_));
  AND4_X1   g345(.A1(new_n537_), .A2(new_n540_), .A3(new_n542_), .A4(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G99gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n539_), .A3(KEYINPUT64), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT7), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n551_), .A2(new_n548_), .A3(new_n539_), .A4(KEYINPUT64), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n537_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  INV_X1    g353(.A(new_n541_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n545_), .A2(KEYINPUT65), .A3(new_n541_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT8), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT8), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n553_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n547_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT73), .B1(new_n532_), .B2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n540_), .A2(new_n537_), .A3(new_n542_), .A4(new_n546_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n563_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n562_), .B1(new_n553_), .B2(new_n559_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT73), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n518_), .A4(new_n520_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(KEYINPUT35), .ZN(new_n574_));
  INV_X1    g373(.A(new_n508_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n564_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n565_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(KEYINPUT35), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(KEYINPUT74), .A3(new_n579_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n569_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n586_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n585_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n596_), .A2(new_n590_), .A3(new_n589_), .A4(new_n583_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n594_), .A2(KEYINPUT37), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n597_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n605_));
  XOR2_X1   g404(.A(G71gat), .B(G78gat), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n564_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT66), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n569_), .A2(new_n608_), .A3(new_n607_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT67), .ZN(new_n613_));
  OAI211_X1 g412(.A(G230gat), .B(G233gat), .C1(new_n611_), .C2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT69), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n569_), .B2(KEYINPUT68), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n612_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G120gat), .B(G148gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n622_), .A2(new_n627_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n602_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n630_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(KEYINPUT13), .A3(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n609_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(new_n493_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT16), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT17), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT17), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n637_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT78), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n637_), .B(KEYINPUT68), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n642_), .B(KEYINPUT77), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n601_), .A2(new_n634_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n531_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n483_), .A3(new_n335_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n594_), .A2(new_n597_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT103), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT104), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n482_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n634_), .A2(new_n530_), .A3(new_n650_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G1gat), .B1(new_n662_), .B2(new_n336_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n653_), .A2(new_n654_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n655_), .A2(new_n663_), .A3(new_n664_), .ZN(G1324gat));
  AND2_X1   g464(.A1(new_n416_), .A2(new_n422_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G8gat), .B1(new_n662_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT39), .ZN(new_n668_));
  INV_X1    g467(.A(new_n666_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n652_), .A2(new_n484_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n662_), .B2(new_n481_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT41), .Z(new_n675_));
  INV_X1    g474(.A(new_n338_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n285_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n652_), .A2(new_n269_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(G1326gat));
  OAI21_X1  g478(.A(G22gat), .B1(new_n662_), .B2(new_n448_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT42), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n448_), .A2(G22gat), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT105), .Z(new_n683_));
  NAND2_X1  g482(.A1(new_n652_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1327gat));
  INV_X1    g484(.A(new_n650_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n657_), .A2(new_n686_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n687_), .A2(new_n482_), .A3(new_n530_), .A4(new_n634_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n335_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n634_), .A2(new_n530_), .A3(new_n686_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n416_), .A2(new_n422_), .A3(new_n451_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n479_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n481_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n666_), .A2(new_n336_), .A3(new_n677_), .A4(new_n448_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n691_), .B1(new_n696_), .B2(new_n601_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT43), .B(new_n600_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n690_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  INV_X1    g501(.A(new_n690_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n482_), .B2(new_n600_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n696_), .A2(new_n691_), .A3(new_n601_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n700_), .B1(new_n706_), .B2(KEYINPUT106), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n690_), .B(KEYINPUT106), .C1(new_n697_), .C2(new_n698_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n702_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT44), .B1(new_n699_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(KEYINPUT107), .A3(new_n708_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n701_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n336_), .A2(new_n496_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n689_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n688_), .A2(new_n494_), .A3(new_n669_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n701_), .A2(new_n666_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n699_), .A2(new_n711_), .ZN(new_n720_));
  AND4_X1   g519(.A1(KEYINPUT107), .A2(new_n720_), .A3(new_n700_), .A4(new_n708_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n712_), .B2(new_n708_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT108), .B(new_n719_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n710_), .A2(new_n713_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT108), .B1(new_n725_), .B2(new_n719_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n718_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT46), .B(new_n718_), .C1(new_n724_), .C2(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n714_), .A2(G43gat), .A3(new_n677_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(G43gat), .ZN(new_n733_));
  INV_X1    g532(.A(new_n688_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n481_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n688_), .B2(new_n479_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n448_), .A2(new_n499_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n714_), .B2(new_n742_), .ZN(G1331gat));
  NAND4_X1  g542(.A1(new_n660_), .A2(new_n530_), .A3(new_n634_), .A4(new_n686_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n336_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n696_), .A2(new_n530_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n747_), .A2(new_n634_), .A3(new_n686_), .A4(new_n600_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n336_), .A2(G57gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1332gat));
  OAI21_X1  g549(.A(G64gat), .B1(new_n744_), .B2(new_n666_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT48), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n666_), .A2(G64gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n748_), .B2(new_n753_), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n744_), .B2(new_n481_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT49), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n481_), .A2(G71gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n748_), .B2(new_n757_), .ZN(G1334gat));
  OAI21_X1  g557(.A(G78gat), .B1(new_n744_), .B2(new_n448_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT50), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n448_), .A2(G78gat), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT110), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n748_), .B2(new_n762_), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n704_), .A2(new_n705_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n634_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n530_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n686_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n543_), .B1(new_n769_), .B2(new_n335_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n746_), .A2(new_n687_), .A3(new_n765_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n336_), .A2(G85gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT111), .ZN(G1336gat));
  AOI21_X1  g573(.A(G92gat), .B1(new_n771_), .B2(new_n669_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT112), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n768_), .A2(new_n544_), .A3(new_n666_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1337gat));
  AOI21_X1  g577(.A(new_n548_), .B1(new_n769_), .B2(new_n677_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n771_), .A2(new_n677_), .A3(new_n538_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n779_), .A2(KEYINPUT113), .A3(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n769_), .A2(new_n479_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G106gat), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT52), .B(new_n539_), .C1(new_n769_), .C2(new_n479_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n771_), .A2(new_n539_), .A3(new_n479_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1339gat));
  NAND2_X1  g590(.A1(new_n651_), .A2(new_n530_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(KEYINPUT54), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(KEYINPUT54), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n621_), .B2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n617_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n620_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n621_), .A2(new_n798_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n620_), .A2(new_n610_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(G230gat), .A3(G233gat), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .A4(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n627_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n627_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n509_), .A2(new_n510_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n513_), .A2(new_n511_), .A3(new_n521_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n527_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n529_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n813_), .B2(new_n812_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n632_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT58), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n809_), .A2(KEYINPUT58), .A3(new_n816_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n601_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n601_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n817_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n815_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT118), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n815_), .B(new_n830_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n807_), .A2(KEYINPUT116), .A3(new_n808_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n804_), .A2(new_n834_), .A3(KEYINPUT56), .A4(new_n627_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n630_), .A2(new_n530_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n832_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n657_), .B1(new_n839_), .B2(KEYINPUT57), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n827_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n838_), .A2(new_n827_), .A3(new_n840_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n822_), .B(new_n825_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n796_), .B1(new_n844_), .B2(new_n650_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n666_), .A2(new_n335_), .A3(new_n448_), .A4(new_n677_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847_), .B2(new_n766_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n846_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n820_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n796_), .B1(new_n851_), .B2(new_n650_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n846_), .A2(KEYINPUT59), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n850_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n650_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n795_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT121), .A3(new_n853_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n849_), .A2(new_n855_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n209_), .B1(new_n766_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n860_), .B2(new_n209_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n848_), .B1(new_n859_), .B2(new_n862_), .ZN(G1340gat));
  NAND4_X1  g662(.A1(new_n849_), .A2(new_n855_), .A3(new_n858_), .A4(new_n634_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G120gat), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT60), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT123), .B1(new_n866_), .B2(G120gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(G120gat), .B1(new_n634_), .B2(new_n866_), .ZN(new_n868_));
  MUX2_X1   g667(.A(new_n867_), .B(KEYINPUT123), .S(new_n868_), .Z(new_n869_));
  NAND2_X1  g668(.A1(new_n847_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n870_), .ZN(G1341gat));
  NAND4_X1  g670(.A1(new_n849_), .A2(new_n855_), .A3(new_n858_), .A4(new_n686_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G127gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n847_), .A2(new_n204_), .A3(new_n686_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  NAND4_X1  g674(.A1(new_n849_), .A2(new_n855_), .A3(new_n858_), .A4(new_n601_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G134gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n847_), .A2(new_n202_), .A3(new_n659_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1343gat));
  NOR2_X1   g678(.A1(new_n845_), .A2(new_n677_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n669_), .A2(new_n336_), .A3(new_n448_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n766_), .A3(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n634_), .A3(new_n881_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g684(.A1(new_n880_), .A2(new_n686_), .A3(new_n881_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1346gat));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n881_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G162gat), .B1(new_n889_), .B2(new_n600_), .ZN(new_n890_));
  INV_X1    g689(.A(G162gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n659_), .A2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n889_), .B2(new_n892_), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n666_), .A2(new_n339_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n479_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n852_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n857_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT22), .B(G169gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n766_), .A3(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n857_), .A2(new_n766_), .A3(new_n896_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n904_), .A2(new_n905_), .A3(G169gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(G169gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n903_), .B1(new_n906_), .B2(new_n907_), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n901_), .A2(new_n634_), .ZN(new_n909_));
  INV_X1    g708(.A(G176gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n845_), .A2(new_n479_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n765_), .A2(new_n895_), .A3(new_n910_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n909_), .A2(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  NOR2_X1   g712(.A1(new_n650_), .A2(new_n261_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n686_), .A3(new_n894_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n901_), .A2(new_n914_), .B1(new_n915_), .B2(new_n252_), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n659_), .A2(new_n251_), .A3(new_n349_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT125), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n901_), .A2(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n600_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n348_), .ZN(G1351gat));
  NOR3_X1   g720(.A1(new_n666_), .A2(new_n335_), .A3(new_n448_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n880_), .A2(new_n766_), .A3(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g723(.A1(new_n880_), .A2(new_n634_), .A3(new_n922_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT126), .B(G204gat), .Z(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1353gat));
  AND2_X1   g726(.A1(new_n844_), .A2(new_n650_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n481_), .B(new_n922_), .C1(new_n928_), .C2(new_n796_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(KEYINPUT127), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(KEYINPUT127), .ZN(new_n932_));
  NAND2_X1  g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n686_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  OR3_X1    g733(.A1(new_n929_), .A2(new_n931_), .A3(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n931_), .B1(new_n929_), .B2(new_n934_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1354gat));
  OAI21_X1  g736(.A(G218gat), .B1(new_n929_), .B2(new_n600_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n659_), .A2(new_n363_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n929_), .B2(new_n939_), .ZN(G1355gat));
endmodule


