//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_;
  NAND2_X1  g000(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(G228gat), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT88), .B(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(G204gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G211gat), .B(G218gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n210_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n212_), .B1(G197gat), .B2(G204gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(KEYINPUT21), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(KEYINPUT89), .B2(new_n211_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n222_), .B(new_n208_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(KEYINPUT90), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G197gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT88), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT88), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G197gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n210_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT89), .B1(new_n229_), .B2(new_n207_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n214_), .A2(KEYINPUT21), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n223_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT90), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n219_), .B1(new_n224_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT84), .B1(new_n238_), .B2(KEYINPUT1), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT84), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(G155gat), .A4(G162gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(KEYINPUT1), .ZN(new_n243_));
  OR2_X1    g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n239_), .A2(new_n242_), .A3(new_n243_), .A4(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G141gat), .B(G148gat), .Z(new_n246_));
  AOI21_X1  g045(.A(new_n237_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n237_), .A3(new_n246_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  OR3_X1    g049(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n252_));
  INV_X1    g051(.A(G141gat), .ZN(new_n253_));
  INV_X1    g052(.A(G148gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT86), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n251_), .B(new_n252_), .C1(new_n255_), .C2(KEYINPUT2), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n255_), .A2(KEYINPUT2), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n238_), .B(new_n244_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n236_), .B1(new_n250_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n206_), .B1(new_n235_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT90), .B1(new_n221_), .B2(new_n223_), .ZN(new_n261_));
  AND4_X1   g060(.A1(KEYINPUT90), .A2(new_n230_), .A3(new_n231_), .A4(new_n223_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n218_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n249_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n258_), .B1(new_n264_), .B2(new_n247_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT29), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n266_), .A3(new_n205_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT91), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G78gat), .B(G106gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n269_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT28), .B1(new_n265_), .B2(KEYINPUT29), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n250_), .A2(new_n275_), .A3(new_n236_), .A4(new_n258_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G22gat), .B(G50gat), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n273_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n268_), .A2(new_n271_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n260_), .A2(new_n267_), .A3(new_n272_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(KEYINPUT91), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n268_), .A2(new_n288_), .A3(new_n271_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n289_), .A2(new_n284_), .A3(new_n280_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n287_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n289_), .A2(new_n284_), .A3(new_n280_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n294_), .A2(KEYINPUT93), .A3(new_n291_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n286_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297_));
  XOR2_X1   g096(.A(G8gat), .B(G36gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G169gat), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(KEYINPUT24), .A3(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n306_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G183gat), .ZN(new_n314_));
  INV_X1    g113(.A(G190gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT23), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(G183gat), .A3(G190gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(KEYINPUT83), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n320_), .A2(new_n317_), .A3(G183gat), .A4(G190gat), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n317_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n316_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n314_), .A2(new_n315_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n311_), .A2(KEYINPUT80), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(G169gat), .A3(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n307_), .A2(KEYINPUT22), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n307_), .A2(KEYINPUT22), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n336_), .B2(new_n308_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n313_), .A2(new_n322_), .B1(new_n328_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT96), .B1(new_n235_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT96), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n263_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n329_), .A2(new_n331_), .A3(new_n309_), .A4(KEYINPUT24), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n306_), .A2(new_n310_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n347_));
  AOI21_X1  g146(.A(G176gat), .B1(new_n333_), .B2(KEYINPUT82), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n332_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n319_), .A2(new_n327_), .A3(new_n321_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n345_), .A2(new_n326_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(new_n218_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT20), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT95), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n355_), .A3(KEYINPUT20), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n343_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT94), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n218_), .B(new_n338_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n361_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n365_), .A2(KEYINPUT20), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT97), .B1(new_n235_), .B2(new_n351_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT97), .ZN(new_n369_));
  INV_X1    g168(.A(new_n351_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n263_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n303_), .B1(new_n363_), .B2(new_n373_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n302_), .B(new_n372_), .C1(new_n357_), .C2(new_n362_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n297_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n362_), .ZN(new_n377_));
  AND4_X1   g176(.A1(new_n377_), .A2(new_n343_), .A3(new_n354_), .A4(new_n356_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n368_), .A2(new_n371_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n235_), .B2(new_n338_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n365_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n302_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n363_), .A2(new_n303_), .A3(new_n373_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT101), .A4(KEYINPUT27), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n376_), .A2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n372_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n297_), .B1(new_n387_), .B2(new_n303_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT101), .B1(new_n388_), .B2(new_n383_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT102), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT27), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT101), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT102), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(new_n376_), .A4(new_n385_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n296_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G71gat), .B(G99gat), .ZN(new_n397_));
  INV_X1    g196(.A(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n351_), .B(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G127gat), .B(G134gat), .Z(new_n401_));
  XOR2_X1   g200(.A(G113gat), .B(G120gat), .Z(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n400_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(G15gat), .Z(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT30), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n404_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n403_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n250_), .A3(new_n258_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n265_), .A2(new_n403_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT4), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n265_), .A2(new_n416_), .A3(new_n403_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n414_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(new_n411_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G85gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT0), .B(G57gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n418_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n410_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n290_), .A2(new_n287_), .A3(new_n292_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT93), .B1(new_n294_), .B2(new_n291_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n432_), .A2(new_n433_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n436_));
  OAI211_X1 g235(.A(KEYINPUT33), .B(new_n425_), .C1(new_n418_), .C2(new_n420_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT99), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n411_), .B1(new_n419_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n438_), .B2(new_n419_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n415_), .A2(new_n411_), .A3(new_n417_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n426_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n443_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI211_X1 g245(.A(new_n446_), .B(new_n372_), .C1(new_n357_), .C2(new_n362_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n379_), .A2(new_n381_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n361_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n343_), .A2(new_n354_), .A3(new_n377_), .A4(new_n356_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n445_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n429_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n434_), .B1(new_n444_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n393_), .A2(new_n376_), .A3(new_n385_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n296_), .A2(new_n429_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n396_), .A2(new_n431_), .B1(new_n456_), .B2(new_n409_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G29gat), .B(G36gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G43gat), .B(G50gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT75), .B(G8gat), .Z(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n460_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n464_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n465_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n460_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n466_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n460_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n472_), .A2(new_n466_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n469_), .B(new_n476_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  NAND3_X1  g284(.A1(new_n478_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n478_), .A2(new_n482_), .A3(KEYINPUT79), .A4(new_n485_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n478_), .A2(new_n482_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n485_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n457_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(G230gat), .A2(G233gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT64), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT6), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR4_X1   g307(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n502_), .B(new_n504_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT66), .B1(new_n516_), .B2(new_n511_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT8), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n515_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n510_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n517_), .ZN(new_n521_));
  INV_X1    g320(.A(G99gat), .ZN(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n507_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT65), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n506_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n525_), .A2(new_n526_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n503_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT6), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT67), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(KEYINPUT67), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(KEYINPUT6), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n503_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n521_), .B1(new_n527_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n520_), .B1(new_n538_), .B2(new_n518_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n542_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT10), .B(G99gat), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n523_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n512_), .A2(KEYINPUT9), .A3(new_n514_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n514_), .A2(KEYINPUT9), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n504_), .A4(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n539_), .A2(new_n546_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT68), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n539_), .A2(new_n554_), .A3(new_n546_), .A4(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n521_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n502_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n534_), .A2(new_n535_), .A3(new_n503_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n503_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n558_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT8), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n557_), .B1(new_n564_), .B2(new_n520_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(new_n546_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n497_), .B1(new_n556_), .B2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n497_), .B1(new_n565_), .B2(new_n546_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT69), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT12), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n539_), .A2(new_n551_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n546_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n574_));
  AOI211_X1 g373(.A(new_n546_), .B(new_n574_), .C1(new_n539_), .C2(new_n551_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n568_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n567_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G120gat), .B(G148gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT71), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n567_), .A2(new_n576_), .A3(new_n582_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(KEYINPUT72), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT34), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n480_), .B1(new_n539_), .B2(new_n551_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n539_), .A2(new_n460_), .A3(new_n551_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT35), .B(new_n596_), .C1(new_n597_), .C2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n480_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n571_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .A4(new_n598_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(KEYINPUT74), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT73), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n600_), .A2(new_n613_), .A3(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n607_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n594_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n618_), .A2(KEYINPUT37), .A3(new_n614_), .A4(new_n612_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n546_), .B(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(new_n481_), .Z(new_n628_));
  AOI211_X1 g427(.A(new_n621_), .B(new_n625_), .C1(new_n628_), .C2(KEYINPUT76), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(KEYINPUT76), .B2(new_n628_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n625_), .B(new_n621_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n628_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n632_), .B2(new_n628_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n630_), .A2(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n593_), .A2(new_n620_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT78), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n496_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G1gat), .A3(new_n429_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n615_), .A2(new_n616_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n457_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n592_), .A2(new_n494_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT103), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n635_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n429_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n640_), .A2(new_n641_), .A3(new_n650_), .ZN(G1324gat));
  AND2_X1   g450(.A1(new_n390_), .A2(new_n395_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n648_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT39), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n461_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n638_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  OAI21_X1  g458(.A(G15gat), .B1(new_n649_), .B2(new_n409_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT105), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n662_), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n638_), .A2(G15gat), .A3(new_n409_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(G1326gat));
  OAI21_X1  g465(.A(G22gat), .B1(new_n649_), .B2(new_n434_), .ZN(new_n667_));
  XOR2_X1   g466(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n434_), .A2(G22gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n638_), .B2(new_n670_), .ZN(G1327gat));
  NAND2_X1  g470(.A1(new_n617_), .A2(new_n619_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n457_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n456_), .A2(new_n409_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n296_), .B(new_n430_), .C1(new_n390_), .C2(new_n395_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n674_), .B(new_n620_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n673_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n646_), .A2(new_n635_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT44), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n682_), .B(new_n679_), .C1(new_n673_), .C2(new_n677_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n681_), .A2(new_n683_), .A3(new_n429_), .ZN(new_n684_));
  INV_X1    g483(.A(G29gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n643_), .A2(new_n635_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n593_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n496_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n429_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n685_), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n684_), .A2(new_n685_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1328gat));
  NAND2_X1  g492(.A1(new_n390_), .A2(new_n395_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT109), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT110), .B1(new_n688_), .B2(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n496_), .A4(new_n687_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n697_), .A2(KEYINPUT45), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT45), .B1(new_n697_), .B2(new_n700_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n681_), .A2(new_n683_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n652_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n694_), .A2(new_n434_), .A3(new_n431_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n456_), .A2(new_n409_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n674_), .B1(new_n709_), .B2(new_n620_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT43), .B(new_n672_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n680_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n682_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n678_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(new_n704_), .A3(new_n652_), .A4(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n703_), .B1(new_n706_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n703_), .B(KEYINPUT46), .C1(new_n706_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NOR3_X1   g520(.A1(new_n681_), .A2(new_n683_), .A3(new_n409_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n410_), .A2(new_n398_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n722_), .A2(new_n398_), .B1(new_n688_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(G1330gat));
  INV_X1    g525(.A(new_n688_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G50gat), .B1(new_n727_), .B2(new_n296_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n296_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n705_), .B2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n457_), .A2(new_n494_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n620_), .A2(new_n635_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n731_), .A2(new_n593_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n689_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n635_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n592_), .A2(new_n494_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n644_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n429_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(new_n739_), .ZN(G1332gat));
  OAI21_X1  g539(.A(G64gat), .B1(new_n738_), .B2(new_n695_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  INV_X1    g543(.A(new_n695_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n733_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n738_), .B2(new_n409_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n733_), .A2(new_n751_), .A3(new_n410_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n738_), .B2(new_n434_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n733_), .A2(new_n756_), .A3(new_n296_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n737_), .A2(new_n635_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n673_), .B2(new_n677_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n429_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n686_), .A2(new_n592_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n731_), .A2(new_n763_), .ZN(new_n764_));
  OR3_X1    g563(.A1(new_n764_), .A2(G85gat), .A3(new_n429_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n761_), .B2(new_n695_), .ZN(new_n767_));
  OR3_X1    g566(.A1(new_n764_), .A2(G92gat), .A3(new_n694_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n761_), .B2(new_n409_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n410_), .A2(new_n547_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n764_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g572(.A(new_n523_), .B1(new_n760_), .B2(new_n296_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT114), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n759_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n296_), .B(new_n777_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n775_), .A3(G106gat), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n434_), .B(new_n759_), .C1(new_n673_), .C2(new_n677_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n782_), .B(KEYINPUT52), .C1(new_n783_), .C2(new_n523_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n778_), .A2(KEYINPUT113), .A3(new_n775_), .A4(G106gat), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n776_), .A2(new_n781_), .A3(new_n784_), .A4(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n731_), .A2(new_n523_), .A3(new_n296_), .A4(new_n763_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  OAI21_X1  g591(.A(new_n469_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n476_), .B1(new_n793_), .B2(KEYINPUT118), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(KEYINPUT118), .B2(new_n793_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n485_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n490_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n573_), .A2(new_n575_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n497_), .B1(new_n800_), .B2(new_n556_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n576_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n568_), .B(KEYINPUT55), .C1(new_n573_), .C2(new_n575_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n801_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n583_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n583_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n494_), .A2(new_n585_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n583_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(KEYINPUT117), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n799_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n643_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n808_), .A2(new_n810_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n585_), .A2(new_n490_), .A3(new_n797_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n672_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(KEYINPUT58), .A3(new_n818_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n816_), .A2(KEYINPUT57), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n799_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n583_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n825_), .A2(new_n813_), .A3(KEYINPUT117), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n806_), .A2(KEYINPUT117), .A3(new_n807_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n812_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n642_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT119), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT119), .B(new_n832_), .C1(new_n815_), .C2(new_n643_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n823_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n736_), .B1(new_n836_), .B2(KEYINPUT120), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n823_), .B(new_n838_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n732_), .A2(new_n495_), .A3(new_n592_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n840_), .B2(KEYINPUT54), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n636_), .A2(new_n842_), .A3(new_n843_), .A4(new_n495_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(KEYINPUT54), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT116), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n848_), .A3(KEYINPUT54), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n837_), .A2(new_n839_), .B1(new_n845_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n396_), .A2(new_n689_), .A3(new_n410_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n845_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n823_), .B1(KEYINPUT57), .B2(new_n816_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n635_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n852_), .A2(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n853_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n494_), .A2(G113gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT123), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT121), .B1(new_n851_), .B2(new_n852_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n836_), .A2(KEYINPUT120), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n635_), .A3(new_n839_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n854_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  INV_X1    g667(.A(new_n852_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n870_), .A3(new_n494_), .ZN(new_n871_));
  INV_X1    g670(.A(G113gat), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(KEYINPUT122), .A3(new_n872_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n863_), .B1(new_n875_), .B2(new_n876_), .ZN(G1340gat));
  AND2_X1   g676(.A1(new_n864_), .A2(new_n870_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n592_), .A2(KEYINPUT60), .ZN(new_n879_));
  MUX2_X1   g678(.A(new_n879_), .B(KEYINPUT60), .S(G120gat), .Z(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n853_), .A2(new_n593_), .A3(new_n859_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G120gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n883_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n881_), .B1(new_n885_), .B2(new_n886_), .ZN(G1341gat));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n878_), .A2(new_n888_), .A3(new_n736_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G127gat), .B1(new_n860_), .B2(new_n635_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1342gat));
  AOI21_X1  g690(.A(new_n852_), .B1(new_n866_), .B2(new_n854_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n620_), .B(new_n859_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G134gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n642_), .A2(G134gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n864_), .A2(new_n870_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT125), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n900_), .A3(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1343gat));
  NOR2_X1   g701(.A1(new_n851_), .A2(new_n410_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n745_), .A2(new_n434_), .A3(new_n429_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n495_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n253_), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n592_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n254_), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n903_), .A2(new_n736_), .A3(new_n904_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT61), .B(G155gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1346gat));
  OAI21_X1  g711(.A(G162gat), .B1(new_n905_), .B2(new_n672_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n642_), .A2(G162gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n905_), .B2(new_n914_), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n695_), .A2(new_n430_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n857_), .A2(new_n434_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n307_), .B1(new_n918_), .B2(new_n494_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n919_), .A2(KEYINPUT62), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n918_), .A2(new_n336_), .A3(new_n494_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(KEYINPUT62), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(G1348gat));
  AOI21_X1  g722(.A(G176gat), .B1(new_n918_), .B2(new_n593_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n851_), .A2(new_n296_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n916_), .A2(G176gat), .A3(new_n593_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n925_), .B2(new_n927_), .ZN(G1349gat));
  NOR3_X1   g727(.A1(new_n917_), .A2(new_n304_), .A3(new_n635_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n925_), .A2(new_n736_), .A3(new_n916_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n314_), .B2(new_n930_), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n917_), .B2(new_n672_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n643_), .A2(new_n305_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n917_), .B2(new_n933_), .ZN(G1351gat));
  NOR2_X1   g733(.A1(new_n695_), .A2(new_n455_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n903_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n495_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n225_), .ZN(G1352gat));
  INV_X1    g737(.A(new_n936_), .ZN(new_n939_));
  XOR2_X1   g738(.A(KEYINPUT126), .B(G204gat), .Z(new_n940_));
  NAND3_X1  g739(.A1(new_n939_), .A2(new_n593_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n210_), .A2(KEYINPUT126), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n936_), .B2(new_n592_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n903_), .A2(new_n736_), .A3(new_n935_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n945_), .A2(new_n946_), .A3(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  XOR2_X1   g748(.A(KEYINPUT127), .B(G218gat), .Z(new_n950_));
  NOR3_X1   g749(.A1(new_n936_), .A2(new_n672_), .A3(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n939_), .A2(new_n643_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n950_), .ZN(G1355gat));
endmodule


