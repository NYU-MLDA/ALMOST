//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(G218gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G211gat), .ZN(new_n204_));
  INV_X1    g003(.A(G211gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G218gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT92), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n210_), .A2(new_n211_), .A3(G204gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(G197gat), .B2(G204gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n208_), .A2(new_n209_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(G204gat), .B1(new_n210_), .B2(new_n211_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G197gat), .A2(G204gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT21), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n204_), .A2(new_n206_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT92), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n217_), .A2(KEYINPUT21), .A3(new_n219_), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n216_), .A2(new_n220_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(G228gat), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT87), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G141gat), .A2(G148gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT89), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT89), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n238_), .B1(new_n248_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n239_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(new_n250_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n236_), .B1(new_n235_), .B2(KEYINPUT1), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n233_), .A2(new_n261_), .A3(new_n234_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n259_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n256_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT29), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n226_), .B(new_n230_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n230_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n268_));
  INV_X1    g067(.A(new_n238_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n246_), .A2(new_n247_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n242_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  NOR4_X1   g073(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(new_n252_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n269_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n234_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT1), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n262_), .A3(new_n237_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n258_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n268_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n211_), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT91), .A2(G197gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n222_), .A2(new_n223_), .B1(new_n287_), .B2(new_n214_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n220_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n225_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n208_), .A2(new_n209_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n288_), .A2(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n267_), .B1(new_n283_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT94), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n266_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n266_), .B2(new_n293_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n202_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n266_), .A2(new_n293_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT94), .ZN(new_n299_));
  INV_X1    g098(.A(new_n202_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n266_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n264_), .A2(new_n304_), .A3(new_n265_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n277_), .A2(new_n282_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n306_), .B2(KEYINPUT29), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G22gat), .B(G50gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n310_), .A2(KEYINPUT95), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n309_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT95), .B1(new_n310_), .B2(new_n311_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n303_), .B2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G8gat), .B(G36gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT18), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT101), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT25), .B(G183gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n329_), .A2(new_n330_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336_));
  INV_X1    g135(.A(G183gat), .ZN(new_n337_));
  INV_X1    g136(.A(G190gat), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n335_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n339_), .B(new_n340_), .C1(G183gat), .C2(G190gat), .ZN(new_n343_));
  AND3_X1   g142(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT22), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT22), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G169gat), .ZN(new_n350_));
  INV_X1    g149(.A(G176gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n343_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n342_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n226_), .B1(new_n328_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(new_n353_), .A3(KEYINPUT101), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n327_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(G169gat), .B1(new_n349_), .B2(KEYINPUT82), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n347_), .A3(KEYINPUT22), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n360_), .A3(new_n351_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n346_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT83), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n364_), .A3(new_n346_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n365_), .A3(new_n343_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n346_), .A2(new_n332_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(G183gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n337_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n370_), .B(new_n371_), .C1(KEYINPUT25), .C2(new_n337_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT26), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n341_), .B(new_n367_), .C1(new_n372_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n366_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n226_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n326_), .B1(new_n357_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n327_), .B1(new_n226_), .B2(new_n354_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n288_), .A2(new_n289_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n290_), .A2(new_n291_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n366_), .A2(new_n380_), .A3(new_n381_), .A4(new_n375_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n325_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n323_), .B1(new_n378_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n323_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n325_), .A2(new_n327_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n377_), .B(new_n387_), .C1(new_n226_), .C2(new_n354_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT96), .B1(new_n383_), .B2(new_n325_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT96), .ZN(new_n390_));
  AOI211_X1 g189(.A(new_n390_), .B(new_n326_), .C1(new_n379_), .C2(new_n382_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n386_), .B(new_n388_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(KEYINPUT27), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT103), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n323_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n392_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n394_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  AOI211_X1 g199(.A(KEYINPUT103), .B(new_n398_), .C1(new_n396_), .C2(new_n392_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n319_), .B(new_n393_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(G15gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n376_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(G43gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n405_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n405_), .A2(new_n411_), .ZN(new_n413_));
  INV_X1    g212(.A(G134gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(G127gat), .ZN(new_n415_));
  INV_X1    g214(.A(G127gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G134gat), .ZN(new_n417_));
  INV_X1    g216(.A(G120gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G113gat), .ZN(new_n419_));
  INV_X1    g218(.A(G113gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G120gat), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n415_), .A2(new_n417_), .A3(new_n419_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n415_), .A2(new_n417_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT31), .Z(new_n426_));
  NAND3_X1  g225(.A1(new_n412_), .A2(new_n413_), .A3(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(KEYINPUT85), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(KEYINPUT85), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI211_X1 g231(.A(KEYINPUT86), .B(new_n426_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n428_), .A2(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G1gat), .B(G29gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G85gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT0), .B(G57gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n425_), .B1(new_n256_), .B2(new_n263_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT97), .B1(new_n423_), .B2(new_n424_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n415_), .A2(new_n417_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n419_), .A2(new_n421_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT97), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n422_), .A3(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n277_), .A2(new_n282_), .A3(new_n440_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n439_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT99), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n439_), .A2(new_n446_), .A3(KEYINPUT99), .A4(new_n447_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n306_), .A2(new_n454_), .A3(new_n425_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n447_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n439_), .A2(new_n446_), .A3(KEYINPUT4), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT98), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT98), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n439_), .A2(new_n446_), .A3(new_n460_), .A4(KEYINPUT4), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n457_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n438_), .B1(new_n453_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n461_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n457_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n438_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n434_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n402_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n438_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n452_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n455_), .A2(new_n447_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n439_), .A2(new_n446_), .A3(new_n456_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n438_), .ZN(new_n479_));
  OAI22_X1  g278(.A1(new_n475_), .A2(new_n462_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT33), .B1(new_n466_), .B2(new_n467_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n482_), .A2(KEYINPUT100), .A3(new_n392_), .A4(new_n396_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT100), .ZN(new_n484_));
  INV_X1    g283(.A(new_n438_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n452_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n473_), .B1(new_n486_), .B2(new_n462_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n477_), .A2(new_n479_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n466_), .A2(new_n452_), .A3(new_n474_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n484_), .B1(new_n490_), .B2(new_n397_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n378_), .B2(new_n384_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n469_), .B(new_n493_), .C1(new_n395_), .C2(new_n492_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n483_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n319_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n318_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n297_), .A2(new_n302_), .A3(new_n312_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n497_), .A2(new_n498_), .A3(new_n469_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(new_n393_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n434_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n472_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT73), .B(G1gat), .ZN(new_n504_));
  INV_X1    g303(.A(G8gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT74), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G8gat), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n510_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G29gat), .B(G36gat), .Z(new_n514_));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n516_), .B(KEYINPUT15), .Z(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n512_), .A3(new_n511_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT78), .Z(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n513_), .B(new_n516_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n521_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n523_), .B(new_n528_), .C1(new_n524_), .C2(new_n521_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n503_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n535_));
  NOR2_X1   g334(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G120gat), .B(G148gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT5), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G176gat), .B(G204gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G85gat), .ZN(new_n543_));
  INV_X1    g342(.A(G92gat), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n543_), .A2(new_n544_), .A3(KEYINPUT9), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G85gat), .B(G92gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(KEYINPUT9), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT10), .B(G99gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n548_), .B1(G106gat), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n546_), .B(KEYINPUT67), .Z(new_n556_));
  OR2_X1    g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557_));
  AND2_X1   g356(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n558_));
  NOR2_X1   g357(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n556_), .B1(new_n553_), .B2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n555_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(KEYINPUT69), .A3(KEYINPUT12), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT68), .B(G71gat), .ZN(new_n567_));
  INV_X1    g366(.A(G78gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G57gat), .B(G64gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(KEYINPUT11), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n573_), .B1(new_n576_), .B2(new_n569_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n579_), .B(new_n555_), .C1(new_n563_), .C2(new_n564_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n566_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n565_), .A2(KEYINPUT69), .A3(KEYINPUT12), .A4(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G230gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT64), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n565_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n578_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n565_), .A2(new_n577_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n542_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n591_), .A3(new_n542_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n537_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n596_), .A2(new_n592_), .A3(new_n535_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n513_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n578_), .ZN(new_n602_));
  XOR2_X1   g401(.A(KEYINPUT69), .B(KEYINPUT75), .Z(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n603_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n605_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n610_), .B(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n602_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n588_), .A2(new_n517_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT35), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI22_X1  g421(.A1(new_n565_), .A2(new_n519_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n618_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT72), .ZN(new_n629_));
  XOR2_X1   g428(.A(G134gat), .B(G162gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n624_), .A2(new_n625_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n626_), .A2(new_n627_), .A3(new_n631_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n631_), .B(KEYINPUT36), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n626_), .B2(new_n632_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n634_), .A2(new_n637_), .A3(KEYINPUT37), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT37), .ZN(new_n639_));
  INV_X1    g438(.A(new_n637_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(new_n633_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n534_), .A2(new_n599_), .A3(new_n616_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n469_), .A3(new_n504_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n634_), .A2(new_n637_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n503_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n613_), .A2(new_n615_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n598_), .A2(new_n653_), .A3(new_n533_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n470_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n650_), .A3(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(new_n393_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n400_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n401_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n646_), .A2(new_n505_), .A3(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n652_), .A2(new_n662_), .A3(new_n654_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n663_), .B(new_n670_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n655_), .B2(new_n502_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT41), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n644_), .A2(G15gat), .A3(new_n502_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n655_), .B2(new_n319_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n319_), .A2(G22gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n644_), .B2(new_n682_), .ZN(G1327gat));
  NAND3_X1  g482(.A1(new_n599_), .A2(new_n532_), .A3(new_n653_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n661_), .A2(new_n499_), .B1(new_n495_), .B2(new_n319_), .ZN(new_n687_));
  OAI22_X1  g486(.A1(new_n687_), .A2(new_n434_), .B1(new_n402_), .B2(new_n471_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(new_n642_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n434_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n686_), .B(new_n642_), .C1(new_n690_), .C2(new_n472_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n685_), .B1(new_n689_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT43), .B1(new_n503_), .B2(new_n643_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n684_), .B1(new_n698_), .B2(new_n691_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT109), .B1(new_n699_), .B2(new_n695_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(KEYINPUT44), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n469_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G29gat), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n653_), .A2(new_n651_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n598_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n534_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n469_), .A2(new_n704_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT110), .Z(new_n709_));
  OAI22_X1  g508(.A1(new_n703_), .A2(new_n704_), .B1(new_n707_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(G36gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n661_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n701_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n707_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n661_), .A2(G36gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n717_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n718_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n719_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n707_), .B2(new_n722_), .ZN(new_n723_));
  AOI22_X1  g522(.A1(new_n720_), .A2(new_n723_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n713_), .B1(new_n716_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n713_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n702_), .A2(new_n662_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n700_), .B2(new_n697_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n727_), .B(new_n724_), .C1(new_n729_), .C2(new_n714_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n726_), .A2(new_n730_), .ZN(G1329gat));
  OAI21_X1  g530(.A(new_n407_), .B1(new_n707_), .B2(new_n502_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT113), .Z(new_n733_));
  NOR2_X1   g532(.A1(new_n502_), .A2(new_n407_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n701_), .A2(new_n702_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n733_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1330gat));
  INV_X1    g540(.A(new_n319_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G50gat), .B1(new_n717_), .B2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n701_), .A2(new_n702_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n742_), .A2(G50gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(new_n651_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n653_), .A2(new_n532_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n688_), .A2(new_n598_), .A3(new_n747_), .A4(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n652_), .A2(KEYINPUT115), .A3(new_n598_), .A4(new_n748_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(G57gat), .A3(new_n469_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n754_), .A2(new_n755_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n503_), .A2(new_n532_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n599_), .A2(new_n653_), .A3(new_n642_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n469_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n756_), .A2(new_n757_), .A3(new_n762_), .ZN(G1332gat));
  OR3_X1    g562(.A1(new_n760_), .A2(G64gat), .A3(new_n661_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n753_), .A2(new_n662_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G64gat), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT48), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  OR3_X1    g568(.A1(new_n760_), .A2(G71gat), .A3(new_n502_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n751_), .A2(new_n752_), .A3(new_n434_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G71gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT117), .ZN(G1334gat));
  NAND3_X1  g575(.A1(new_n761_), .A2(new_n568_), .A3(new_n742_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n753_), .A2(new_n742_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G78gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n705_), .A2(new_n599_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n758_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n543_), .A3(new_n469_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n698_), .A2(new_n691_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n599_), .A2(new_n616_), .A3(new_n532_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n789_), .A2(new_n469_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n790_), .B2(new_n543_), .ZN(G1336gat));
  NAND3_X1  g590(.A1(new_n785_), .A2(new_n544_), .A3(new_n662_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n789_), .A2(new_n662_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n544_), .ZN(G1337gat));
  NAND2_X1  g593(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n502_), .A2(new_n549_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n784_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n789_), .A2(new_n434_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(G99gat), .ZN(new_n799_));
  NOR2_X1   g598(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1338gat));
  OR3_X1    g600(.A1(new_n784_), .A2(G106gat), .A3(new_n319_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n742_), .A3(new_n788_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(G106gat), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n803_), .B2(G106gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n616_), .A2(new_n809_), .A3(new_n533_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n642_), .A2(new_n598_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT119), .B1(new_n653_), .B2(new_n532_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .A4(new_n814_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n522_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n518_), .A2(new_n520_), .A3(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n529_), .C1(new_n524_), .C2(new_n819_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n531_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n587_), .A2(KEYINPUT55), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n583_), .A2(new_n825_), .A3(new_n586_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n583_), .A2(new_n586_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT56), .B(new_n541_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  INV_X1    g629(.A(new_n583_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n824_), .A2(new_n826_), .B1(new_n831_), .B2(new_n585_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n832_), .B2(new_n542_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n532_), .A2(new_n835_), .A3(new_n594_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n532_), .B2(new_n594_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n823_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT122), .B1(new_n839_), .B2(new_n651_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT57), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n596_), .A2(new_n822_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT58), .B1(new_n834_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n643_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n834_), .A2(KEYINPUT58), .A3(new_n842_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT122), .B(new_n847_), .C1(new_n839_), .C2(new_n651_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n841_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n818_), .B1(new_n849_), .B2(new_n653_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n402_), .A2(new_n470_), .A3(new_n502_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT123), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n851_), .A2(new_n420_), .A3(new_n532_), .A4(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  INV_X1    g654(.A(new_n853_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n850_), .B2(new_n856_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n840_), .A2(KEYINPUT57), .B1(new_n844_), .B2(new_n845_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n616_), .B1(new_n858_), .B2(new_n848_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT59), .B(new_n853_), .C1(new_n859_), .C2(new_n818_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n533_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n854_), .B1(new_n861_), .B2(new_n420_), .ZN(G1340gat));
  NOR2_X1   g661(.A1(new_n850_), .A2(new_n856_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n418_), .B1(new_n599_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n863_), .B(new_n864_), .C1(KEYINPUT60), .C2(new_n418_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n599_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n418_), .ZN(G1341gat));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n416_), .A3(new_n616_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n653_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n416_), .ZN(G1342gat));
  NAND3_X1  g669(.A1(new_n863_), .A2(new_n414_), .A3(new_n651_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n643_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n414_), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n434_), .A2(new_n319_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n661_), .A2(new_n874_), .A3(new_n469_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT124), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n851_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877_), .B2(new_n533_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n876_), .ZN(new_n879_));
  OR4_X1    g678(.A1(G141gat), .A2(new_n850_), .A3(new_n533_), .A4(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1344gat));
  OAI21_X1  g680(.A(G148gat), .B1(new_n877_), .B2(new_n599_), .ZN(new_n882_));
  OR4_X1    g681(.A1(G148gat), .A2(new_n850_), .A3(new_n599_), .A4(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1345gat));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n877_), .B2(new_n653_), .ZN(new_n886_));
  OR4_X1    g685(.A1(new_n653_), .A2(new_n850_), .A3(new_n879_), .A4(new_n885_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1346gat));
  INV_X1    g687(.A(G162gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n651_), .A2(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n850_), .A2(new_n643_), .A3(new_n879_), .ZN(new_n891_));
  OAI22_X1  g690(.A1(new_n877_), .A2(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1347gat));
  NAND3_X1  g691(.A1(new_n434_), .A2(new_n319_), .A3(new_n470_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n661_), .A2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n532_), .B(new_n894_), .C1(new_n859_), .C2(new_n818_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G169gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n894_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n850_), .A2(new_n899_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n900_), .A2(new_n348_), .A3(new_n350_), .A4(new_n532_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n895_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n900_), .B2(new_n598_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n850_), .A2(new_n351_), .A3(new_n599_), .A4(new_n899_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1349gat));
  NOR4_X1   g705(.A1(new_n850_), .A2(new_n329_), .A3(new_n653_), .A4(new_n899_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n900_), .A2(new_n616_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n337_), .B2(new_n908_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n900_), .A2(new_n330_), .A3(new_n651_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n850_), .A2(new_n643_), .A3(new_n899_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n338_), .B2(new_n911_), .ZN(G1351gat));
  NAND3_X1  g711(.A1(new_n662_), .A2(new_n470_), .A3(new_n874_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n850_), .A2(new_n533_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  NOR3_X1   g715(.A1(new_n850_), .A2(new_n599_), .A3(new_n913_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n285_), .ZN(G1353gat));
  NOR2_X1   g717(.A1(new_n850_), .A2(new_n913_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n653_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT125), .Z(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT126), .Z(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n919_), .A2(new_n920_), .A3(new_n924_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1354gat));
  AOI21_X1  g727(.A(G218gat), .B1(new_n919_), .B2(new_n651_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n642_), .A2(G218gat), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n930_), .B(KEYINPUT127), .Z(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n919_), .B2(new_n931_), .ZN(G1355gat));
endmodule


