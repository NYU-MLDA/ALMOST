//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n212_), .B(KEYINPUT87), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n219_), .B(new_n220_), .C1(G183gat), .C2(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n206_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n217_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT21), .B1(new_n226_), .B2(KEYINPUT83), .ZN(new_n227_));
  XOR2_X1   g026(.A(G197gat), .B(G204gat), .Z(new_n228_));
  OAI211_X1 g027(.A(new_n227_), .B(new_n228_), .C1(KEYINPUT21), .C2(new_n226_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT21), .B(new_n230_), .C1(new_n226_), .C2(KEYINPUT83), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT20), .B(new_n204_), .C1(new_n225_), .C2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT78), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n222_), .A2(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n206_), .B1(new_n236_), .B2(KEYINPUT78), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n221_), .B(new_n212_), .C1(new_n235_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n216_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n232_), .A3(KEYINPUT88), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n233_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n239_), .A2(new_n232_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT20), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n225_), .B2(new_n232_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n204_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G8gat), .B(G36gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT18), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G64gat), .B(G92gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n250_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n242_), .A2(new_n243_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n232_), .A2(KEYINPUT84), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n229_), .A2(new_n263_), .A3(new_n231_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n261_), .B(KEYINPUT20), .C1(new_n265_), .C2(new_n225_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n203_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n246_), .A2(new_n248_), .A3(new_n204_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT93), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n254_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n255_), .A2(KEYINPUT27), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n260_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G78gat), .B(G106gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT86), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT2), .ZN(new_n279_));
  OR2_X1    g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT3), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(KEYINPUT2), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(KEYINPUT3), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT81), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(G155gat), .A3(G162gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n284_), .B(new_n289_), .C1(G155gat), .C2(G162gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n280_), .A2(new_n276_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(KEYINPUT1), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(G155gat), .B2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n289_), .A2(KEYINPUT1), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n291_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT29), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n265_), .ZN(new_n298_));
  INV_X1    g097(.A(G228gat), .ZN(new_n299_));
  INV_X1    g098(.A(G233gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(KEYINPUT85), .A3(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n297_), .B(new_n232_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n275_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n296_), .A2(KEYINPUT29), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT28), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(KEYINPUT28), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G22gat), .B(G50gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n306_), .A2(new_n275_), .A3(new_n307_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n309_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n315_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n306_), .A2(new_n275_), .A3(new_n307_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(new_n308_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n272_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G134gat), .Z(new_n328_));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND3_X1  g129(.A1(new_n296_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT91), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n296_), .A2(new_n330_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n330_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(new_n290_), .A3(new_n295_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(KEYINPUT4), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT90), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n335_), .A2(new_n340_), .A3(KEYINPUT4), .A4(new_n337_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n334_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n335_), .A2(new_n337_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(G225gat), .B2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G1gat), .B(G29gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  INV_X1    g152(.A(new_n351_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(KEYINPUT94), .B(new_n354_), .C1(new_n342_), .C2(new_n345_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT79), .B(G43gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(G15gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G71gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n362_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT31), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT80), .B1(new_n336_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n369_), .B2(new_n336_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G99gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n368_), .B(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n326_), .A2(new_n359_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n320_), .A2(new_n324_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n244_), .A2(new_n249_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n378_), .B2(new_n376_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n352_), .A2(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n255_), .A2(KEYINPUT89), .A3(new_n257_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT89), .B1(new_n255_), .B2(new_n257_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n343_), .A2(KEYINPUT33), .A3(new_n346_), .A4(new_n351_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n339_), .A2(new_n341_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n332_), .A3(new_n331_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n333_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n388_), .B(new_n354_), .C1(new_n344_), .C2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n382_), .A2(new_n385_), .A3(new_n386_), .A4(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n375_), .A2(new_n380_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n272_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n373_), .B1(new_n393_), .B2(new_n375_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT96), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n320_), .A2(new_n324_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n272_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n358_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n375_), .A2(new_n380_), .A3(new_n391_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .A4(new_n373_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n374_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G8gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT72), .ZN(new_n405_));
  INV_X1    g204(.A(G22gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n364_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G15gat), .A2(G22gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G1gat), .A2(G8gat), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n407_), .A2(new_n408_), .B1(KEYINPUT14), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n405_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G29gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n414_), .B2(new_n411_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n411_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n414_), .B(KEYINPUT15), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G229gat), .A2(G233gat), .ZN(new_n423_));
  MUX2_X1   g222(.A(new_n418_), .B(new_n422_), .S(new_n423_), .Z(new_n424_));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(G113gat), .B(G141gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT76), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G169gat), .B(G197gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n424_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n403_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G85gat), .ZN(new_n437_));
  INV_X1    g236(.A(G92gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n439_), .B(new_n440_), .C1(new_n441_), .C2(KEYINPUT65), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(KEYINPUT65), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT68), .B1(new_n444_), .B2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n441_), .A2(KEYINPUT65), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n439_), .A2(new_n440_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n441_), .A2(KEYINPUT65), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n448_), .A2(new_n453_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G85gat), .B(G92gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n464_));
  INV_X1    g263(.A(G99gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n446_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI211_X1 g267(.A(KEYINPUT8), .B(new_n463_), .C1(new_n468_), .C2(new_n453_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n453_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n463_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n455_), .B(new_n462_), .C1(new_n469_), .C2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n450_), .A2(new_n452_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n466_), .A2(new_n467_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n472_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n482_), .A2(KEYINPUT69), .A3(new_n455_), .A4(new_n462_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n420_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n459_), .A2(new_n460_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n486_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G232gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT71), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n488_), .A2(new_n414_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n485_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n494_), .A2(new_n489_), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  XNOR2_X1  g297(.A(G190gat), .B(G218gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G134gat), .B(G162gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(KEYINPUT36), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n501_), .B(KEYINPUT36), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(KEYINPUT37), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(KEYINPUT37), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G127gat), .B(G155gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G183gat), .B(G211gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT17), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(KEYINPUT17), .ZN(new_n515_));
  XOR2_X1   g314(.A(G71gat), .B(G78gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(KEYINPUT11), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n517_), .B2(KEYINPUT11), .ZN(new_n520_));
  INV_X1    g319(.A(G64gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(G57gat), .ZN(new_n522_));
  INV_X1    g321(.A(G57gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(G64gat), .ZN(new_n524_));
  AND4_X1   g323(.A1(new_n519_), .A2(new_n522_), .A3(new_n524_), .A4(KEYINPUT11), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n518_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n524_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT11), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT66), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n519_), .A3(KEYINPUT11), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n528_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .A4(new_n516_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(new_n419_), .ZN(new_n536_));
  MUX2_X1   g335(.A(new_n514_), .B(new_n515_), .S(new_n536_), .Z(new_n537_));
  XOR2_X1   g336(.A(new_n537_), .B(KEYINPUT74), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n508_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n526_), .A2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT12), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n476_), .B2(new_n483_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT12), .B1(new_n487_), .B2(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT64), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n487_), .B2(new_n540_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT67), .B1(new_n487_), .B2(new_n540_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n482_), .A2(new_n533_), .A3(new_n549_), .A4(new_n486_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n488_), .B2(new_n533_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n545_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n547_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G120gat), .B(G148gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G176gat), .B(G204gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n559_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n539_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n436_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(G1gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n359_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT97), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT38), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT98), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n572_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT100), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n505_), .B(KEYINPUT99), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n403_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n435_), .A2(new_n566_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n538_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n584_), .B2(new_n358_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n574_), .A2(new_n576_), .A3(new_n585_), .ZN(G1324gat));
  OAI21_X1  g385(.A(G8gat), .B1(new_n584_), .B2(new_n397_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT39), .ZN(new_n588_));
  INV_X1    g387(.A(G8gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n568_), .A2(new_n589_), .A3(new_n272_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g391(.A(new_n584_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n373_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n364_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n568_), .A2(new_n364_), .A3(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(G1326gat));
  OAI21_X1  g399(.A(G22gat), .B1(new_n584_), .B2(new_n375_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n568_), .A2(new_n406_), .A3(new_n396_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1327gat));
  NOR3_X1   g404(.A1(new_n566_), .A2(new_n538_), .A3(new_n505_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n436_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(G29gat), .B1(new_n608_), .B2(new_n359_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n403_), .A2(KEYINPUT43), .A3(new_n508_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n395_), .A2(new_n402_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n374_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT103), .ZN(new_n616_));
  INV_X1    g415(.A(new_n508_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n403_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n616_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n612_), .B1(new_n620_), .B2(KEYINPUT43), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n403_), .B2(new_n618_), .ZN(new_n622_));
  AOI211_X1 g421(.A(KEYINPUT103), .B(new_n374_), .C1(new_n395_), .C2(new_n402_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n612_), .B(KEYINPUT43), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n611_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n581_), .A2(new_n538_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT44), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n622_), .B2(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT104), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n610_), .B1(new_n632_), .B2(new_n624_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n627_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n628_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n359_), .A2(G29gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n609_), .B1(new_n636_), .B2(new_n637_), .ZN(G1328gat));
  NAND3_X1  g437(.A1(new_n628_), .A2(new_n635_), .A3(new_n272_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G36gat), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n397_), .A2(KEYINPUT106), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n397_), .A2(KEYINPUT106), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n607_), .A2(G36gat), .A3(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT45), .Z(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n640_), .A2(KEYINPUT46), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1329gat));
  NAND4_X1  g450(.A1(new_n628_), .A2(new_n635_), .A3(G43gat), .A4(new_n594_), .ZN(new_n652_));
  INV_X1    g451(.A(G43gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n607_), .B2(new_n373_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g455(.A(G50gat), .B1(new_n608_), .B2(new_n396_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n396_), .A2(G50gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n636_), .B2(new_n658_), .ZN(G1331gat));
  NAND2_X1  g458(.A1(new_n615_), .A2(new_n435_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT108), .ZN(new_n661_));
  INV_X1    g460(.A(new_n566_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n539_), .A2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT107), .Z(new_n664_));
  AND2_X1   g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n523_), .A3(new_n359_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n662_), .A2(new_n434_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n579_), .A2(new_n538_), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G57gat), .B1(new_n668_), .B2(new_n358_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1332gat));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n521_), .A3(new_n643_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G64gat), .B1(new_n668_), .B2(new_n644_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT48), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1333gat));
  OAI21_X1  g473(.A(G71gat), .B1(new_n668_), .B2(new_n373_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT109), .Z(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT49), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT49), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n665_), .A2(new_n366_), .A3(new_n594_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(G1334gat));
  INV_X1    g479(.A(G78gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n665_), .A2(new_n681_), .A3(new_n396_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G78gat), .B1(new_n668_), .B2(new_n375_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT50), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1335gat));
  NOR3_X1   g484(.A1(new_n662_), .A2(new_n505_), .A3(new_n538_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n661_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT110), .B1(new_n661_), .B2(new_n686_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n437_), .A3(new_n359_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n667_), .A2(new_n582_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT112), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n626_), .B2(KEYINPUT111), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n633_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n696_), .A2(new_n358_), .A3(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n692_), .B1(new_n699_), .B2(new_n437_), .ZN(G1336gat));
  NAND3_X1  g499(.A1(new_n691_), .A2(new_n438_), .A3(new_n272_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n696_), .A2(new_n644_), .A3(new_n698_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(new_n438_), .ZN(G1337gat));
  AND3_X1   g502(.A1(new_n594_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n691_), .A2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n696_), .A2(new_n373_), .A3(new_n698_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n465_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT51), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n705_), .B(new_n709_), .C1(new_n706_), .C2(new_n465_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1338gat));
  NAND2_X1  g510(.A1(new_n695_), .A2(new_n396_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G106gat), .B1(new_n633_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT114), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT114), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(G106gat), .C1(new_n633_), .C2(new_n712_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n714_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n713_), .A2(KEYINPUT114), .A3(new_n717_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n689_), .A2(new_n690_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n375_), .A2(G106gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT53), .B1(new_n719_), .B2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n691_), .A2(new_n722_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .A4(new_n720_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1339gat));
  NAND2_X1  g529(.A1(new_n567_), .A2(new_n435_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT54), .Z(new_n732_));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n733_));
  INV_X1    g532(.A(new_n541_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n484_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n543_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n551_), .A3(new_n736_), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n553_), .A2(new_n737_), .B1(new_n547_), .B2(KEYINPUT55), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n547_), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT115), .ZN(new_n740_));
  INV_X1    g539(.A(new_n546_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n736_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n739_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT116), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT115), .B1(new_n547_), .B2(KEYINPUT55), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n740_), .A3(new_n743_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n738_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n559_), .B1(new_n746_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n733_), .B1(new_n752_), .B2(KEYINPUT56), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT56), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n749_), .A2(new_n750_), .A3(new_n738_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n750_), .B1(new_n749_), .B2(new_n738_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n558_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(KEYINPUT117), .A3(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n754_), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n418_), .B1(G229gat), .B2(G233gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n422_), .A2(new_n423_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n430_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n554_), .B2(new_n559_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n760_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n760_), .A2(KEYINPUT58), .A3(new_n765_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n617_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n434_), .A2(new_n561_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n757_), .A2(new_n758_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n754_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n764_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT57), .B(new_n505_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n505_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n770_), .A2(new_n775_), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n732_), .B1(new_n582_), .B2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n326_), .A2(new_n358_), .A3(new_n373_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n784_));
  INV_X1    g583(.A(new_n775_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n770_), .A2(new_n778_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(KEYINPUT118), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n770_), .A2(new_n788_), .A3(new_n778_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n538_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n732_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n781_), .A2(new_n784_), .ZN(new_n792_));
  OAI22_X1  g591(.A1(new_n783_), .A2(new_n784_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G113gat), .B1(new_n793_), .B2(new_n435_), .ZN(new_n794_));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n795_), .A3(new_n434_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1340gat));
  OAI21_X1  g596(.A(G120gat), .B1(new_n793_), .B2(new_n662_), .ZN(new_n798_));
  INV_X1    g597(.A(G120gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n662_), .B2(KEYINPUT60), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n783_), .B(new_n800_), .C1(KEYINPUT60), .C2(new_n799_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n801_), .ZN(G1341gat));
  OAI21_X1  g601(.A(G127gat), .B1(new_n793_), .B2(new_n582_), .ZN(new_n803_));
  INV_X1    g602(.A(G127gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n783_), .A2(new_n804_), .A3(new_n538_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1342gat));
  NOR3_X1   g605(.A1(new_n780_), .A2(new_n577_), .A3(new_n782_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n807_), .A2(KEYINPUT119), .A3(G134gat), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(G134gat), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(G134gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n508_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI221_X1 g611(.A(new_n812_), .B1(new_n791_), .B2(new_n792_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT119), .B1(new_n807_), .B2(G134gat), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n808_), .A2(new_n813_), .A3(new_n814_), .ZN(G1343gat));
  NAND2_X1  g614(.A1(new_n396_), .A2(new_n373_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n780_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n643_), .A2(new_n358_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n435_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT121), .B(G141gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1344gat));
  INV_X1    g621(.A(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n566_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n538_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  OR3_X1    g627(.A1(new_n819_), .A2(G162gat), .A3(new_n577_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G162gat), .B1(new_n819_), .B2(new_n508_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1347gat));
  NOR2_X1   g630(.A1(new_n359_), .A2(new_n373_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n643_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n396_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n791_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n205_), .B1(new_n836_), .B2(new_n434_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT122), .A3(KEYINPUT62), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n434_), .A2(new_n222_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT123), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n838_), .B(new_n841_), .C1(new_n837_), .C2(new_n842_), .ZN(G1348gat));
  AOI21_X1  g642(.A(G176gat), .B1(new_n836_), .B2(new_n566_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n780_), .A2(new_n396_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n833_), .A2(new_n206_), .A3(new_n662_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1349gat));
  NAND4_X1  g646(.A1(new_n845_), .A2(new_n832_), .A3(new_n538_), .A4(new_n643_), .ZN(new_n848_));
  INV_X1    g647(.A(G183gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n582_), .A2(new_n209_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n848_), .A2(new_n849_), .B1(new_n836_), .B2(new_n850_), .ZN(G1350gat));
  NAND3_X1  g650(.A1(new_n836_), .A2(new_n210_), .A3(new_n578_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n617_), .B(new_n834_), .C1(new_n790_), .C2(new_n732_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(new_n854_), .A3(G190gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n853_), .B2(G190gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n852_), .B(KEYINPUT125), .C1(new_n855_), .C2(new_n856_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1351gat));
  NOR2_X1   g660(.A1(new_n644_), .A2(new_n359_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n817_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G197gat), .B1(new_n864_), .B2(new_n434_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n817_), .A2(G197gat), .A3(new_n434_), .A4(new_n862_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(KEYINPUT126), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(KEYINPUT126), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n864_), .A2(new_n566_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g670(.A(KEYINPUT63), .B(G211gat), .C1(new_n864_), .C2(new_n538_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT63), .B(G211gat), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n863_), .A2(new_n582_), .A3(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1354gat));
  AOI21_X1  g674(.A(G218gat), .B1(new_n864_), .B2(new_n578_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n617_), .A2(G218gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT127), .Z(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n864_), .B2(new_n878_), .ZN(G1355gat));
endmodule


