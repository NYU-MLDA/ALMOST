//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G71gat), .B(G78gat), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n206_), .A3(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G127gat), .B(G155gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(G211gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT16), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT17), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT75), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G231gat), .ZN(new_n217_));
  INV_X1    g016(.A(G233gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G8gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G22gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT73), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT73), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G22gat), .ZN(new_n227_));
  INV_X1    g026(.A(G15gat), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT74), .ZN(new_n232_));
  XOR2_X1   g031(.A(G1gat), .B(G8gat), .Z(new_n233_));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n234_), .B(new_n223_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n233_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n215_), .A2(new_n219_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n221_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n238_), .B1(new_n221_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n209_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n221_), .A2(new_n239_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n209_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n221_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n213_), .A2(KEYINPUT17), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n242_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G141gat), .A2(G148gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT2), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n254_));
  OR3_X1    g053(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT86), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G155gat), .B(G162gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  INV_X1    g060(.A(G141gat), .ZN(new_n262_));
  INV_X1    g061(.A(G148gat), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n261_), .A2(KEYINPUT1), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n252_), .C1(KEYINPUT1), .C2(new_n258_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G113gat), .B(G120gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n260_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT4), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(new_n275_), .C1(KEYINPUT4), .C2(new_n271_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n274_), .A3(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G57gat), .B(G85gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G29gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n276_), .A2(new_n277_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT87), .B(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(G197gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n293_), .B(KEYINPUT21), .C1(new_n292_), .C2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(G197gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(G197gat), .B2(new_n294_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n295_), .B(new_n296_), .C1(new_n298_), .C2(KEYINPUT21), .ZN(new_n299_));
  INV_X1    g098(.A(new_n296_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(KEYINPUT21), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT23), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT22), .B(G169gat), .Z(new_n308_));
  OAI211_X1 g107(.A(new_n306_), .B(new_n307_), .C1(G176gat), .C2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT26), .B(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(G183gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT25), .B(G183gat), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n310_), .B(new_n313_), .C1(new_n314_), .C2(new_n311_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(KEYINPUT24), .A3(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT78), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n305_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT79), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n315_), .A2(KEYINPUT78), .A3(new_n318_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n321_), .A2(new_n326_), .A3(new_n327_), .A4(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n303_), .A2(new_n309_), .A3(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n324_), .A2(KEYINPUT92), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n324_), .A2(KEYINPUT92), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n310_), .A2(new_n314_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n318_), .A4(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n309_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n302_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n331_), .A2(new_n337_), .A3(KEYINPUT20), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT20), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n330_), .A2(new_n309_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(new_n302_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n303_), .A2(new_n309_), .A3(new_n335_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n349_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n290_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n331_), .A2(new_n337_), .A3(KEYINPUT20), .A4(new_n341_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT98), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n346_), .A2(new_n347_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n343_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n355_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n365_), .A2(new_n366_), .B1(new_n355_), .B2(new_n350_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT27), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n360_), .A2(KEYINPUT98), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n360_), .A2(KEYINPUT98), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n357_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n368_), .B1(new_n372_), .B2(KEYINPUT99), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n359_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(G50gat), .B1(new_n266_), .B2(KEYINPUT29), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT28), .B(G22gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  INV_X1    g176(.A(G50gat), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n260_), .A2(new_n377_), .A3(new_n378_), .A4(new_n265_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n375_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n376_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n303_), .B1(new_n266_), .B2(KEYINPUT29), .ZN(new_n385_));
  INV_X1    g184(.A(G228gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n218_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n385_), .A2(new_n388_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n390_), .A2(KEYINPUT90), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n266_), .A2(KEYINPUT29), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n302_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n387_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n393_), .B1(new_n396_), .B2(new_n389_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n383_), .B(new_n384_), .C1(new_n392_), .C2(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n384_), .B(KEYINPUT88), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n389_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n383_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n399_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n382_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n380_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n405_), .A2(new_n407_), .A3(KEYINPUT89), .A4(new_n401_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n398_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G227gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G43gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(G15gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT80), .B(KEYINPUT82), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n413_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n330_), .A2(new_n419_), .A3(new_n309_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n345_), .A2(KEYINPUT30), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT84), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(KEYINPUT84), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(new_n421_), .A3(new_n420_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT83), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT85), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n426_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n269_), .B(KEYINPUT31), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT85), .B(new_n435_), .C1(new_n425_), .C2(new_n427_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n409_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n409_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n288_), .B(new_n374_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n350_), .B2(KEYINPUT97), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n364_), .A3(new_n362_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n349_), .B2(KEYINPUT97), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n288_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n271_), .A2(new_n275_), .A3(new_n272_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n283_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT96), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n273_), .B(new_n274_), .C1(KEYINPUT4), .C2(new_n271_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(KEYINPUT96), .A3(new_n283_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n276_), .A2(new_n277_), .A3(new_n285_), .A4(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n356_), .A2(new_n452_), .A3(new_n455_), .A4(new_n358_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n286_), .A2(new_n453_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n409_), .B(new_n440_), .C1(new_n445_), .C2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n251_), .B1(new_n439_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G169gat), .B(G197gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n232_), .A2(new_n235_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n233_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT71), .B(G43gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G29gat), .ZN(new_n470_));
  INV_X1    g269(.A(G36gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G29gat), .A2(G36gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n378_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n378_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n469_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G50gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n467_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n481_), .B1(new_n467_), .B2(new_n482_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G229gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(new_n218_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT15), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n481_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n477_), .A2(KEYINPUT15), .A3(new_n480_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(new_n467_), .A3(new_n482_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n475_), .A2(new_n469_), .A3(new_n476_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n468_), .B1(new_n479_), .B2(new_n474_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n488_), .B(KEYINPUT76), .Z(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n464_), .B1(new_n490_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n464_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n501_), .B(new_n504_), .C1(new_n486_), .C2(new_n489_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G204gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT5), .B(G176gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT66), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n516_));
  INV_X1    g315(.A(G99gat), .ZN(new_n517_));
  INV_X1    g316(.A(G106gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n512_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT65), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT6), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n523_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n523_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n515_), .B(new_n521_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G85gat), .B(G92gat), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT8), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n519_), .A2(new_n512_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n526_), .A2(KEYINPUT6), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n524_), .A2(KEYINPUT65), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n522_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n523_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n534_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n531_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n533_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT10), .B(G99gat), .Z(new_n542_));
  AOI22_X1  g341(.A1(KEYINPUT9), .A2(new_n531_), .B1(new_n542_), .B2(new_n518_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n538_), .ZN(new_n544_));
  INV_X1    g343(.A(G85gat), .ZN(new_n545_));
  INV_X1    g344(.A(G92gat), .ZN(new_n546_));
  OR3_X1    g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT9), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n532_), .A2(new_n541_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n532_), .A2(new_n541_), .A3(new_n548_), .A4(KEYINPUT67), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n246_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n549_), .A2(new_n550_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n552_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n209_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT64), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n246_), .A2(new_n549_), .A3(KEYINPUT12), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n555_), .A2(new_n558_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n560_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n553_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n246_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n511_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n566_), .A3(new_n511_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(KEYINPUT13), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n562_), .A2(new_n566_), .A3(new_n511_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n572_), .B2(new_n567_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n461_), .A2(new_n506_), .A3(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n498_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n494_), .A2(new_n549_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n581_), .A2(new_n582_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n577_), .A2(new_n583_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n481_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n584_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n582_), .B(new_n581_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT72), .ZN(new_n591_));
  XOR2_X1   g390(.A(G190gat), .B(G218gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT36), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT72), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n590_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n576_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n202_), .B1(new_n605_), .B2(new_n287_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT101), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608_));
  INV_X1    g407(.A(new_n595_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n601_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n603_), .B2(new_n608_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n576_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n202_), .A3(new_n287_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n607_), .A2(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(new_n374_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n222_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n605_), .A2(new_n618_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(G8gat), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n621_), .A2(KEYINPUT39), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(KEYINPUT39), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(new_n440_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n228_), .B1(new_n605_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT41), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n614_), .A2(new_n228_), .A3(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1326gat));
  INV_X1    g430(.A(new_n409_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n224_), .B1(new_n605_), .B2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT42), .Z(new_n634_));
  NOR2_X1   g433(.A1(new_n409_), .A2(G22gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT102), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n614_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(G1327gat));
  NAND2_X1  g437(.A1(new_n439_), .A2(new_n460_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n506_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n574_), .A2(new_n640_), .A3(new_n250_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n639_), .A2(new_n604_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT104), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n603_), .B1(new_n439_), .B2(new_n460_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n641_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n287_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n641_), .B(KEYINPUT103), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n639_), .B2(new_n613_), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT43), .B(new_n612_), .C1(new_n439_), .C2(new_n460_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT44), .B(new_n649_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n288_), .A2(new_n470_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n648_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n618_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n647_), .A2(new_n662_), .A3(new_n471_), .A4(new_n618_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n643_), .A2(new_n471_), .A3(new_n618_), .A4(new_n646_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT105), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n663_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n664_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n661_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  OAI221_X1 g471(.A(new_n661_), .B1(new_n670_), .B2(KEYINPUT46), .C1(new_n667_), .C2(new_n668_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  INV_X1    g473(.A(G43gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n647_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n440_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n655_), .A2(G43gat), .A3(new_n627_), .A4(new_n656_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT107), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(KEYINPUT107), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT47), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n683_), .B(new_n677_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1330gat));
  NAND2_X1  g484(.A1(new_n657_), .A2(new_n632_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n657_), .A2(KEYINPUT108), .A3(new_n632_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(G50gat), .A3(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n647_), .A2(new_n378_), .A3(new_n632_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n575_), .A2(new_n506_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n461_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n603_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n696_), .A2(G57gat), .A3(new_n287_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n694_), .A2(new_n612_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n287_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1332gat));
  NOR2_X1   g499(.A1(new_n374_), .A2(G64gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n618_), .A3(new_n603_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G64gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT109), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(G64gat), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n706_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n707_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n703_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT111), .B(new_n703_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n698_), .A2(new_n717_), .A3(new_n627_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n696_), .B2(new_n627_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1334gat));
  OAI21_X1  g522(.A(G78gat), .B1(new_n695_), .B2(new_n409_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n698_), .A2(new_n726_), .A3(new_n632_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1335gat));
  NAND2_X1  g527(.A1(new_n693_), .A2(new_n251_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n603_), .B(new_n729_), .C1(new_n439_), .C2(new_n460_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G85gat), .B1(new_n730_), .B2(new_n287_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n651_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n639_), .A2(new_n650_), .A3(new_n613_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n288_), .A2(new_n545_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1336gat));
  AOI21_X1  g535(.A(G92gat), .B1(new_n730_), .B2(new_n618_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n374_), .A2(new_n546_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n734_), .B2(new_n738_), .ZN(G1337gat));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n542_), .A3(new_n627_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT113), .Z(new_n741_));
  AOI21_X1  g540(.A(new_n517_), .B1(new_n734_), .B2(new_n627_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n743_), .B(new_n744_), .Z(G1338gat));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n409_), .B(new_n729_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n747_), .B2(new_n518_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n734_), .A2(new_n632_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n750_), .A3(KEYINPUT52), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n730_), .A2(new_n518_), .A3(new_n632_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n746_), .B(new_n753_), .C1(new_n747_), .C2(new_n518_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT53), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n751_), .A2(new_n757_), .A3(new_n752_), .A4(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1339gat));
  NOR2_X1   g558(.A1(new_n251_), .A2(new_n506_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n612_), .A2(new_n760_), .A3(new_n575_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n761_), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT116), .B1(new_n761_), .B2(KEYINPUT54), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n500_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n495_), .A2(new_n499_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n464_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n499_), .B2(new_n483_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT117), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n500_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n464_), .A4(new_n767_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n774_), .A2(KEYINPUT118), .A3(new_n505_), .A4(new_n569_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n505_), .A3(new_n773_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n572_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n555_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n563_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n562_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n562_), .A2(KEYINPUT55), .ZN(new_n784_));
  AND4_X1   g583(.A1(KEYINPUT56), .A2(new_n783_), .A3(new_n784_), .A4(new_n510_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n511_), .B1(new_n782_), .B2(new_n562_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n784_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n779_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n779_), .B(KEYINPUT58), .C1(new_n785_), .C2(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n613_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n506_), .A2(new_n569_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n786_), .A2(new_n784_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n784_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n777_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT57), .B(new_n603_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n603_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n790_), .A2(KEYINPUT119), .A3(new_n613_), .A4(new_n791_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n794_), .A2(new_n802_), .A3(new_n805_), .A4(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n765_), .B1(new_n807_), .B2(new_n251_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n618_), .A2(new_n288_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n437_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n506_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT59), .B1(new_n808_), .B2(new_n810_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n808_), .C2(new_n810_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n805_), .A2(new_n792_), .A3(new_n802_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n765_), .B1(new_n251_), .B2(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n819_), .A2(KEYINPUT59), .A3(new_n810_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT121), .B1(new_n817_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n823_), .B(new_n820_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n506_), .A2(G113gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n812_), .B1(new_n825_), .B2(new_n826_), .ZN(G1340gat));
  NOR2_X1   g626(.A1(new_n575_), .A2(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n811_), .B1(KEYINPUT60), .B2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n817_), .A2(new_n574_), .A3(new_n821_), .A4(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(KEYINPUT60), .B2(new_n829_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n811_), .B2(new_n250_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n250_), .A2(G127gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n825_), .B2(new_n834_), .ZN(G1342gat));
  AOI21_X1  g634(.A(G134gat), .B1(new_n811_), .B2(new_n604_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n613_), .A2(G134gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n825_), .B2(new_n837_), .ZN(G1343gat));
  NOR3_X1   g637(.A1(new_n808_), .A2(new_n409_), .A3(new_n627_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n809_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n640_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n262_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n575_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n263_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n840_), .A2(new_n251_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  INV_X1    g646(.A(new_n840_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n848_), .A2(G162gat), .A3(new_n613_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G162gat), .B1(new_n848_), .B2(new_n604_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1347gat));
  NOR2_X1   g650(.A1(new_n374_), .A2(new_n287_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n627_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n640_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT122), .Z(new_n855_));
  NOR3_X1   g654(.A1(new_n855_), .A2(new_n819_), .A3(new_n632_), .ZN(new_n856_));
  INV_X1    g655(.A(G169gat), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n856_), .A2(new_n857_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n859_), .B(new_n863_), .C1(KEYINPUT62), .C2(new_n858_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n818_), .A2(new_n251_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n437_), .B(new_n852_), .C1(new_n865_), .C2(new_n765_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT124), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n867_), .A2(new_n640_), .A3(new_n308_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(G1348gat));
  INV_X1    g668(.A(new_n867_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G176gat), .B1(new_n870_), .B2(new_n574_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n808_), .A2(new_n632_), .ZN(new_n872_));
  INV_X1    g671(.A(G176gat), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n853_), .A2(new_n873_), .A3(new_n575_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n872_), .B2(new_n874_), .ZN(G1349gat));
  NOR2_X1   g674(.A1(new_n853_), .A2(new_n251_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G183gat), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n251_), .A2(new_n314_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n870_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n867_), .B2(new_n612_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n604_), .A2(new_n310_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT125), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n867_), .B2(new_n882_), .ZN(G1351gat));
  AND2_X1   g682(.A1(new_n839_), .A2(new_n852_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n506_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n574_), .ZN(new_n887_));
  MUX2_X1   g686(.A(new_n291_), .B(G204gat), .S(new_n887_), .Z(G1353gat));
  NAND2_X1  g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n250_), .A3(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n890_), .B(new_n893_), .Z(G1354gat));
  AOI21_X1  g693(.A(G218gat), .B1(new_n884_), .B2(new_n604_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n613_), .A2(G218gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n884_), .B2(new_n896_), .ZN(G1355gat));
endmodule


