//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G1gat), .B(G8gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT76), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G1gat), .A2(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT14), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n204_), .A2(KEYINPUT76), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n204_), .A2(KEYINPUT76), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n211_), .A2(new_n208_), .A3(new_n206_), .A4(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G29gat), .B(G36gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n217_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT77), .B1(new_n218_), .B2(new_n219_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n203_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n202_), .B(KEYINPUT78), .Z(new_n225_));
  AND2_X1   g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n217_), .B(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n213_), .A3(new_n210_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G141gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G169gat), .B(G197gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n232_), .B(new_n233_), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT79), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n224_), .A2(new_n237_), .A3(new_n230_), .A4(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n235_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G15gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT87), .B(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G71gat), .B(G99gat), .Z(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT80), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT83), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT83), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT23), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n257_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263_));
  INV_X1    g062(.A(new_n257_), .ZN(new_n264_));
  OAI22_X1  g063(.A1(new_n262_), .A2(new_n263_), .B1(KEYINPUT23), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n266_), .A2(KEYINPUT84), .A3(new_n257_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n256_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT85), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(new_n263_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT84), .B1(new_n266_), .B2(new_n257_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n270_), .B(new_n271_), .C1(KEYINPUT23), .C2(new_n264_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n256_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n255_), .B1(G169gat), .B2(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT81), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT25), .B(G183gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT81), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n275_), .A2(new_n251_), .A3(new_n281_), .A4(new_n253_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT82), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n277_), .A2(new_n285_), .A3(new_n280_), .A4(new_n282_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n269_), .A2(new_n274_), .A3(new_n284_), .A4(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n290_), .B1(new_n264_), .B2(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n259_), .A2(new_n261_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n264_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n266_), .A2(new_n290_), .A3(new_n257_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n289_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n287_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n249_), .B1(new_n300_), .B2(KEYINPUT88), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G134gat), .Z(new_n303_));
  XOR2_X1   g102(.A(G113gat), .B(G120gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n300_), .A2(KEYINPUT88), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n298_), .B(KEYINPUT30), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n302_), .B(new_n307_), .C1(new_n312_), .C2(new_n248_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n307_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n248_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(new_n301_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n320_), .B2(KEYINPUT1), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n321_), .B2(KEYINPUT90), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n323_), .B(new_n318_), .C1(new_n320_), .C2(KEYINPUT1), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(KEYINPUT3), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n326_), .B(KEYINPUT2), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n320_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(new_n318_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT29), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n325_), .A2(new_n329_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT91), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT96), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(KEYINPUT96), .A3(new_n347_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT97), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n345_), .A2(new_n350_), .A3(KEYINPUT97), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n343_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n344_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n348_), .A2(KEYINPUT95), .A3(new_n344_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n362_));
  INV_X1    g161(.A(new_n348_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(KEYINPUT21), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n348_), .A2(KEYINPUT94), .A3(new_n344_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n360_), .B(new_n361_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n356_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n369_), .A2(G228gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(G228gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT93), .Z(new_n373_));
  NAND4_X1  g172(.A1(new_n339_), .A2(new_n342_), .A3(new_n367_), .A4(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n360_), .A2(new_n361_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n364_), .A2(new_n365_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n375_), .A2(new_n376_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n378_));
  NOR2_X1   g177(.A1(new_n340_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n372_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT99), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n340_), .A2(new_n341_), .ZN(new_n385_));
  XOR2_X1   g184(.A(G22gat), .B(G50gat), .Z(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT28), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n385_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n383_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n382_), .B1(new_n374_), .B2(new_n380_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT100), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT100), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n374_), .A2(new_n380_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n381_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n395_), .B2(new_n383_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n389_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT100), .B1(new_n390_), .B2(new_n391_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n393_), .A3(new_n383_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n384_), .A4(new_n388_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n305_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n337_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n340_), .A2(new_n305_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(KEYINPUT103), .Z(new_n407_));
  OR2_X1    g206(.A1(new_n403_), .A2(KEYINPUT4), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT4), .ZN(new_n409_));
  INV_X1    g208(.A(new_n405_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G29gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(G85gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT0), .B(G57gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n406_), .A2(KEYINPUT103), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n406_), .A2(KEYINPUT103), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n418_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n377_), .B1(new_n287_), .B2(new_n297_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT19), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n275_), .A2(KEYINPUT101), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n275_), .A2(KEYINPUT101), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n427_), .A2(new_n253_), .A3(new_n251_), .A4(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n278_), .A2(new_n279_), .B1(new_n255_), .B2(new_n250_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n292_), .A2(new_n264_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n432_), .A2(KEYINPUT84), .B1(new_n258_), .B2(new_n257_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n296_), .B1(new_n433_), .B2(new_n270_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n289_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n426_), .B1(new_n436_), .B2(new_n367_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n423_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT102), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n436_), .B2(new_n367_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n298_), .B2(new_n367_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n439_), .A2(new_n440_), .B1(new_n425_), .B2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT18), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G64gat), .B(G92gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  AOI21_X1  g246(.A(new_n438_), .B1(new_n298_), .B2(new_n367_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n437_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT102), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n447_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n367_), .B1(new_n436_), .B2(KEYINPUT105), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(KEYINPUT105), .B2(new_n436_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n426_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n442_), .A2(new_n425_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n453_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n458_), .A3(KEYINPUT27), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n401_), .A2(new_n422_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n448_), .A2(new_n440_), .A3(new_n449_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n442_), .A2(new_n425_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n439_), .A2(new_n440_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n453_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n447_), .B1(new_n443_), .B2(new_n451_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n461_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT106), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n453_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n452_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(KEYINPUT106), .A3(new_n461_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n460_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n417_), .A2(new_n421_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n447_), .A2(KEYINPUT32), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n443_), .A2(new_n476_), .A3(new_n451_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n456_), .A2(new_n457_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n475_), .B(new_n477_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n408_), .A2(new_n409_), .A3(new_n405_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n403_), .A2(new_n404_), .A3(new_n410_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT104), .A3(new_n416_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT104), .B1(new_n481_), .B2(new_n416_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n421_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n421_), .A2(new_n486_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n487_), .A2(new_n471_), .A3(new_n452_), .A4(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n401_), .B1(new_n479_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n317_), .B1(new_n474_), .B2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n317_), .A2(new_n475_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n470_), .A2(new_n473_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n401_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .A4(new_n459_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n242_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G127gat), .B(G155gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT16), .ZN(new_n499_));
  XOR2_X1   g298(.A(G183gat), .B(G211gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(G231gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n214_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G71gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G71gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(G78gat), .ZN(new_n509_));
  INV_X1    g308(.A(G78gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G57gat), .ZN(new_n513_));
  INV_X1    g312(.A(G57gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(G64gat), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT11), .B1(new_n513_), .B2(new_n515_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n509_), .B(new_n511_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n519_));
  INV_X1    g318(.A(new_n511_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n510_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI211_X1 g323(.A(new_n497_), .B(new_n501_), .C1(new_n503_), .C2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n524_), .B2(new_n503_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n501_), .B(new_n497_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n503_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(KEYINPUT69), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n522_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n532_), .B2(new_n528_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G85gat), .B(G92gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n551_), .B1(G99gat), .B2(G106gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n550_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT67), .B(new_n547_), .C1(new_n555_), .C2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT8), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n551_), .A2(G99gat), .A3(G106gat), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n563_), .A2(new_n564_), .B1(new_n549_), .B2(new_n548_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT67), .B1(new_n566_), .B2(new_n547_), .ZN(new_n567_));
  AOI21_X1  g366(.A(G92gat), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n568_));
  NOR2_X1   g367(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n571_), .A2(KEYINPUT64), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(KEYINPUT64), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n570_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(G106gat), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n577_), .A2(new_n578_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n574_), .A2(new_n579_), .A3(KEYINPUT65), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT65), .B1(new_n574_), .B2(new_n579_), .ZN(new_n581_));
  OAI22_X1  g380(.A1(new_n562_), .A2(new_n567_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n547_), .B1(new_n555_), .B2(new_n560_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT67), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT8), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n545_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n584_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(KEYINPUT8), .A3(new_n561_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n574_), .A2(new_n579_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT65), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n574_), .A2(new_n579_), .A3(KEYINPUT65), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n595_), .A3(KEYINPUT70), .A4(new_n586_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n228_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT74), .B1(new_n542_), .B2(new_n543_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n590_), .A2(new_n595_), .A3(new_n217_), .A4(new_n586_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n544_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n600_), .B(KEYINPUT73), .ZN(new_n605_));
  INV_X1    g404(.A(new_n544_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n603_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n604_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n539_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT37), .B1(new_n608_), .B2(KEYINPUT75), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n603_), .A2(new_n607_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n604_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n603_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n539_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n535_), .B1(new_n612_), .B2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n558_), .A2(new_n559_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n546_), .B1(new_n623_), .B2(new_n565_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n585_), .B1(new_n624_), .B2(KEYINPUT67), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n625_), .A2(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n586_), .A3(new_n532_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n518_), .A2(new_n522_), .A3(new_n530_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n530_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT71), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n532_), .B1(new_n626_), .B2(new_n586_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(KEYINPUT12), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT12), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n524_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n588_), .A2(new_n596_), .A3(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n631_), .A2(KEYINPUT71), .A3(new_n639_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n638_), .A2(new_n627_), .A3(new_n641_), .A4(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n635_), .B1(new_n643_), .B2(new_n634_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT5), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n646_), .B(new_n647_), .Z(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n590_), .A2(new_n586_), .A3(new_n595_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n636_), .B(KEYINPUT12), .C1(new_n650_), .C2(new_n630_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT71), .B1(new_n631_), .B2(new_n639_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n641_), .A2(new_n627_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n633_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n648_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n635_), .A3(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n649_), .A2(KEYINPUT13), .A3(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT13), .B1(new_n649_), .B2(new_n657_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n622_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n496_), .A2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n662_), .A2(G1gat), .A3(new_n422_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT107), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT38), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n610_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n660_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n667_), .A2(new_n242_), .A3(new_n535_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n669_), .B2(new_n422_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(KEYINPUT38), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n665_), .A2(new_n670_), .A3(new_n671_), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n493_), .A2(new_n459_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n666_), .A2(new_n673_), .A3(new_n668_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(KEYINPUT108), .A3(G8gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT108), .B1(new_n674_), .B2(G8gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n676_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(KEYINPUT109), .A2(KEYINPUT39), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n673_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n662_), .A2(G8gat), .A3(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n681_), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n679_), .A2(new_n681_), .A3(new_n683_), .A4(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n669_), .B2(new_n317_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n662_), .A2(G15gat), .A3(new_n317_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n669_), .B2(new_n494_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n494_), .A2(G22gat), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT112), .Z(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n662_), .B2(new_n699_), .ZN(G1327gat));
  NAND4_X1  g499(.A1(new_n496_), .A2(new_n660_), .A3(new_n535_), .A4(new_n610_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n701_), .A2(G29gat), .A3(new_n422_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n612_), .A2(new_n621_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n313_), .A2(new_n316_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n401_), .A2(new_n422_), .A3(new_n459_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT106), .B1(new_n472_), .B2(new_n461_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n469_), .B(KEYINPUT27), .C1(new_n471_), .C2(new_n452_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n479_), .A2(new_n489_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n494_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n705_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n494_), .B(new_n459_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n705_), .A2(new_n422_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n704_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT43), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n491_), .A2(new_n495_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n704_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n535_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n667_), .A2(new_n242_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT44), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  INV_X1    g524(.A(new_n723_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n725_), .B(new_n726_), .C1(new_n717_), .C2(new_n720_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n475_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G29gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n728_), .B2(new_n475_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n702_), .B1(new_n731_), .B2(new_n732_), .ZN(G1328gat));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT115), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT116), .Z(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G36gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n728_), .B2(new_n673_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n673_), .A2(KEYINPUT114), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n673_), .A2(KEYINPUT114), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n738_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n701_), .A2(new_n743_), .A3(KEYINPUT45), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT45), .B1(new_n701_), .B2(new_n743_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n737_), .B1(new_n739_), .B2(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n724_), .A2(new_n727_), .A3(new_n682_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n736_), .B(new_n746_), .C1(new_n749_), .C2(new_n738_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1329gat));
  INV_X1    g550(.A(G43gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n317_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n728_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n701_), .B2(new_n317_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(KEYINPUT47), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT47), .B1(new_n754_), .B2(new_n755_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1330gat));
  INV_X1    g557(.A(G50gat), .ZN(new_n759_));
  NOR4_X1   g558(.A1(new_n724_), .A2(new_n727_), .A3(new_n759_), .A4(new_n494_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n701_), .B2(new_n494_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT117), .B1(new_n760_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n728_), .A2(G50gat), .A3(new_n401_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n761_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(G1331gat));
  AOI21_X1  g566(.A(new_n241_), .B1(new_n491_), .B2(new_n495_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n768_), .A2(new_n667_), .A3(new_n622_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n514_), .A3(new_n475_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n666_), .A2(new_n242_), .A3(new_n667_), .A4(new_n722_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G57gat), .B1(new_n771_), .B2(new_n422_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1332gat));
  INV_X1    g572(.A(new_n742_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G64gat), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT48), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n512_), .A3(new_n742_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n771_), .B2(new_n317_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT49), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n769_), .A2(new_n504_), .A3(new_n705_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1334gat));
  OAI21_X1  g581(.A(G78gat), .B1(new_n771_), .B2(new_n494_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT50), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n401_), .A2(new_n510_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n769_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n784_), .A2(new_n787_), .ZN(G1335gat));
  INV_X1    g587(.A(new_n610_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n660_), .A2(new_n722_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n768_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(G85gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n475_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n721_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n667_), .A2(new_n242_), .A3(new_n535_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n795_), .A2(new_n422_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n794_), .B1(new_n797_), .B2(new_n793_), .ZN(G1336gat));
  INV_X1    g597(.A(G92gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n799_), .A3(new_n673_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n795_), .A2(new_n774_), .A3(new_n796_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n799_), .ZN(G1337gat));
  NAND2_X1  g601(.A1(new_n705_), .A2(new_n577_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n791_), .A2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT119), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n795_), .A2(new_n317_), .A3(new_n796_), .ZN(new_n806_));
  INV_X1    g605(.A(G99gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g608(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n796_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n719_), .B1(new_n718_), .B2(new_n704_), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT43), .B(new_n703_), .C1(new_n491_), .C2(new_n495_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n401_), .B(new_n812_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(G106gat), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(G106gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(KEYINPUT120), .A3(new_n819_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n792_), .A2(new_n578_), .A3(new_n401_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n811_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n818_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT52), .A3(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(new_n822_), .A3(new_n823_), .A4(new_n810_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n829_), .ZN(G1339gat));
  NAND2_X1  g629(.A1(new_n241_), .A2(new_n657_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n643_), .B2(new_n634_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n643_), .A2(new_n634_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n653_), .A2(new_n654_), .A3(KEYINPUT55), .A4(new_n633_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n648_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n633_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n655_), .B1(new_n841_), .B2(new_n832_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n836_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT56), .A3(new_n648_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n831_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n225_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n225_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n234_), .B1(new_n229_), .B2(new_n847_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n236_), .A2(new_n238_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n649_), .A2(new_n657_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n789_), .B1(new_n845_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n789_), .C1(new_n845_), .C2(new_n851_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n849_), .A2(new_n657_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n648_), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n839_), .B(new_n656_), .C1(new_n842_), .C2(new_n836_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n856_), .B(KEYINPUT58), .C1(new_n857_), .C2(new_n858_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n704_), .A3(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n854_), .A2(new_n855_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n535_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n703_), .A2(new_n660_), .A3(new_n242_), .A4(new_n722_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT122), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n622_), .A2(new_n868_), .A3(new_n242_), .A4(new_n660_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n867_), .A2(KEYINPUT54), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT54), .B1(new_n867_), .B2(new_n869_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n317_), .B1(new_n865_), .B2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n713_), .A2(new_n422_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n241_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n873_), .A2(KEYINPUT59), .A3(new_n874_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n242_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n882_), .B2(new_n877_), .ZN(G1340gat));
  INV_X1    g682(.A(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n660_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n876_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n884_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n660_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n884_), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n875_), .B2(new_n535_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n892_), .B(new_n889_), .C1(new_n875_), .C2(new_n535_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n880_), .A2(new_n881_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n535_), .A2(new_n889_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n891_), .A2(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n876_), .A2(new_n897_), .A3(new_n610_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n703_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n705_), .A2(new_n494_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n742_), .A2(new_n422_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n703_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n853_), .A2(new_n852_), .B1(new_n903_), .B2(new_n862_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n722_), .B1(new_n904_), .B2(new_n855_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n867_), .A2(new_n869_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n867_), .A2(KEYINPUT54), .A3(new_n869_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n901_), .B(new_n902_), .C1(new_n905_), .C2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n241_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n667_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g715(.A(KEYINPUT124), .B1(new_n911_), .B2(new_n535_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n901_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n865_), .B2(new_n872_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n722_), .A4(new_n902_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n917_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n917_), .B2(new_n921_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1346gat));
  AOI21_X1  g724(.A(G162gat), .B1(new_n912_), .B2(new_n610_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n704_), .A2(G162gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT125), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n912_), .B2(new_n928_), .ZN(G1347gat));
  INV_X1    g728(.A(KEYINPUT22), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n742_), .A2(new_n422_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n401_), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n873_), .A2(new_n930_), .A3(new_n241_), .A4(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(G169gat), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n933_), .A2(KEYINPUT62), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(KEYINPUT62), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n873_), .A2(new_n937_), .A3(new_n241_), .A4(new_n932_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n938_), .A2(G169gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n936_), .B2(new_n939_), .ZN(G1348gat));
  NAND2_X1  g739(.A1(new_n873_), .A2(new_n932_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(new_n660_), .ZN(new_n942_));
  INV_X1    g741(.A(G176gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1349gat));
  INV_X1    g743(.A(new_n941_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G183gat), .B1(new_n945_), .B2(new_n722_), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n941_), .A2(new_n278_), .A3(new_n535_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n941_), .B2(new_n703_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n610_), .A2(new_n279_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n941_), .B2(new_n950_), .ZN(G1351gat));
  INV_X1    g750(.A(new_n931_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n901_), .B(new_n952_), .C1(new_n905_), .C2(new_n910_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n865_), .A2(new_n872_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n955_), .A2(new_n956_), .A3(new_n901_), .A4(new_n952_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n954_), .A2(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958_), .B2(new_n241_), .ZN(new_n959_));
  INV_X1    g758(.A(G197gat), .ZN(new_n960_));
  AOI211_X1 g759(.A(new_n960_), .B(new_n242_), .C1(new_n954_), .C2(new_n957_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n961_), .ZN(G1352gat));
  NOR2_X1   g761(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n956_), .B1(new_n919_), .B2(new_n952_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n667_), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n967_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n958_), .A2(new_n667_), .A3(new_n966_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(G1353gat));
  NOR2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  INV_X1    g770(.A(new_n971_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n535_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n972_), .B1(new_n958_), .B2(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(new_n973_), .ZN(new_n975_));
  AOI211_X1 g774(.A(new_n971_), .B(new_n975_), .C1(new_n954_), .C2(new_n957_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1354gat));
  INV_X1    g776(.A(G218gat), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n958_), .A2(new_n978_), .A3(new_n610_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n703_), .B1(new_n954_), .B2(new_n957_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n978_), .B2(new_n980_), .ZN(G1355gat));
endmodule


