//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT9), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT64), .A3(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n212_), .C1(new_n209_), .C2(new_n208_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT64), .B1(new_n208_), .B2(new_n209_), .ZN(new_n214_));
  OAI221_X1 g013(.A(new_n206_), .B1(G106gat), .B2(new_n207_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n216_), .B(new_n217_), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n206_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n212_), .A2(new_n208_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n204_), .B(new_n215_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G232gat), .A2(G233gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT34), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT35), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(KEYINPUT35), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT68), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT70), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n215_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT67), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n236_), .B(new_n215_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G190gat), .B(G218gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G134gat), .B(G162gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT36), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n228_), .B1(new_n238_), .B2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n234_), .A2(KEYINPUT69), .A3(new_n235_), .A4(new_n237_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n230_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n239_), .B(new_n243_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n242_), .B(KEYINPUT36), .Z(new_n250_));
  AOI21_X1  g049(.A(new_n248_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n239_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n234_), .A2(new_n237_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G57gat), .B(G64gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G71gat), .B(G78gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(KEYINPUT11), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(KEYINPUT11), .B2(new_n257_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n257_), .A2(KEYINPUT11), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT12), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n256_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G230gat), .A2(G233gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n233_), .A2(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n233_), .A2(new_n264_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT12), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n269_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n267_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT66), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n277_), .A3(new_n274_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n272_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G120gat), .B(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT5), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G176gat), .B(G204gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n283_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n272_), .A2(new_n276_), .A3(new_n278_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT13), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n204_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n235_), .B2(new_n296_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G229gat), .A2(G233gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n289_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n204_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n296_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n304_), .A3(KEYINPUT77), .ZN(new_n305_));
  OR3_X1    g104(.A1(new_n297_), .A2(KEYINPUT77), .A3(new_n204_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n301_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(KEYINPUT78), .B2(new_n308_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G113gat), .B(G141gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G169gat), .B(G197gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n310_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n288_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G183gat), .B(G211gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT73), .ZN(new_n317_));
  XOR2_X1   g116(.A(G127gat), .B(G155gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT72), .B(KEYINPUT16), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT17), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G231gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n296_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(new_n263_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n321_), .A2(new_n322_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n323_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT75), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n328_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT74), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n315_), .A2(KEYINPUT98), .A3(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT98), .B1(new_n315_), .B2(new_n333_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n255_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT82), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT1), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n339_), .B(new_n340_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n341_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n348_), .A2(new_n337_), .A3(new_n338_), .A4(KEYINPUT83), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n350_));
  OAI22_X1  g149(.A1(new_n350_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n340_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  OAI22_X1  g153(.A1(new_n340_), .A2(new_n352_), .B1(new_n348_), .B2(KEYINPUT83), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n347_), .B(new_n343_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n345_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n345_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(KEYINPUT4), .A3(new_n363_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n369_), .A3(new_n361_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n365_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT0), .B(G57gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  OR3_X1    g174(.A1(new_n367_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n371_), .B2(new_n367_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n379_));
  INV_X1    g178(.A(G204gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(G197gat), .ZN(new_n381_));
  INV_X1    g180(.A(G197gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n380_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(G197gat), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G211gat), .B(G218gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT21), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n386_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(G197gat), .B2(G204gat), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n394_), .A2(KEYINPUT85), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT85), .B1(new_n394_), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n384_), .A2(new_n388_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n390_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n393_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT23), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n404_), .A2(KEYINPUT80), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(G183gat), .A3(G190gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT80), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G183gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT25), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT25), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G183gat), .ZN(new_n413_));
  INV_X1    g212(.A(G190gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT26), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT26), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G190gat), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n411_), .A2(new_n413_), .A3(new_n415_), .A4(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G169gat), .A2(G176gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT24), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n418_), .A2(new_n422_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n409_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G176gat), .ZN(new_n428_));
  INV_X1    g227(.A(G169gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT22), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT22), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G169gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n428_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n421_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n404_), .A2(new_n407_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n410_), .A2(new_n414_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n427_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n402_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n389_), .A2(new_n392_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n400_), .A2(new_n390_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449_));
  AND2_X1   g248(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n450_), .A2(new_n451_), .A3(G197gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT21), .B1(new_n382_), .B2(new_n380_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n394_), .A2(KEYINPUT85), .A3(new_n395_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n447_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n442_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n430_), .A2(new_n432_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n440_), .B1(new_n459_), .B2(new_n428_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n438_), .A2(new_n439_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n461_), .A2(new_n420_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n418_), .A2(new_n425_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n458_), .A2(new_n460_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n446_), .A2(new_n465_), .A3(KEYINPUT20), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G226gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT19), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n457_), .A2(new_n464_), .A3(KEYINPUT92), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n458_), .A2(new_n460_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n462_), .A2(new_n463_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n402_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n468_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT20), .B(new_n477_), .C1(new_n402_), .C2(new_n445_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n469_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT18), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  AND2_X1   g282(.A1(new_n483_), .A2(KEYINPUT32), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n378_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT93), .B(KEYINPUT20), .Z(new_n486_));
  AOI22_X1  g285(.A1(new_n409_), .A2(new_n426_), .B1(new_n436_), .B2(new_n443_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n457_), .B2(new_n487_), .ZN(new_n488_));
  OAI22_X1  g287(.A1(new_n470_), .A2(new_n475_), .B1(new_n488_), .B2(KEYINPUT94), .ZN(new_n489_));
  INV_X1    g288(.A(new_n486_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n402_), .B2(new_n445_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n468_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT95), .B1(new_n466_), .B2(new_n468_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n498_), .B(new_n468_), .C1(new_n489_), .C2(new_n493_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n497_), .A2(new_n499_), .A3(new_n484_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT33), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n377_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n377_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n483_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n466_), .A2(new_n468_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT92), .B1(new_n457_), .B2(new_n464_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n402_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n478_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n469_), .B(new_n483_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n375_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n368_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n485_), .A2(new_n500_), .B1(new_n504_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G228gat), .A2(G233gat), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n402_), .B2(KEYINPUT88), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n357_), .A2(KEYINPUT29), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n402_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n520_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n522_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT89), .B1(new_n528_), .B2(new_n523_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n530_));
  AOI211_X1 g329(.A(new_n530_), .B(new_n524_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n527_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G22gat), .B(G50gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n357_), .A2(KEYINPUT29), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n534_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n537_), .A3(new_n533_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n526_), .B2(new_n525_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n528_), .A2(new_n523_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n525_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n532_), .A2(new_n544_), .B1(new_n546_), .B2(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n516_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT27), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n510_), .A2(new_n549_), .A3(new_n511_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n491_), .A2(new_n492_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n488_), .A2(KEYINPUT94), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n477_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n499_), .B(new_n505_), .C1(new_n554_), .C2(new_n495_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n497_), .A2(KEYINPUT96), .A3(new_n505_), .A4(new_n499_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n511_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n551_), .B1(new_n559_), .B2(KEYINPUT27), .ZN(new_n560_));
  INV_X1    g359(.A(new_n527_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n529_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n531_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n544_), .A4(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n546_), .A2(new_n543_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n378_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n548_), .B1(new_n560_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n464_), .B(KEYINPUT30), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G227gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(G15gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G71gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(G99gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n570_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n360_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT81), .B(G43gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT31), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n569_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n559_), .A2(KEYINPUT27), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n566_), .B1(new_n586_), .B2(new_n550_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n378_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n336_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G1gat), .B1(new_n591_), .B2(new_n567_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n253_), .B2(KEYINPUT71), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n254_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n249_), .B(new_n253_), .C1(KEYINPUT71), .C2(new_n594_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n333_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n288_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n314_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n601_), .B2(new_n600_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(new_n590_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT97), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n590_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n567_), .A2(G1gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n593_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n610_), .B2(new_n593_), .ZN(new_n613_));
  OAI221_X1 g412(.A(new_n592_), .B1(new_n593_), .B2(new_n610_), .C1(new_n612_), .C2(new_n613_), .ZN(G1324gat));
  NAND4_X1  g413(.A1(new_n605_), .A2(new_n292_), .A3(new_n560_), .A4(new_n608_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n336_), .A2(new_n590_), .ZN(new_n616_));
  AOI211_X1 g415(.A(KEYINPUT39), .B(new_n292_), .C1(new_n616_), .C2(new_n560_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n560_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(G8gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n615_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n621_), .B(new_n623_), .ZN(G1325gat));
  NAND3_X1  g423(.A1(new_n604_), .A2(new_n572_), .A3(new_n583_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n616_), .A2(new_n583_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n626_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(new_n626_), .B2(G15gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT101), .ZN(G1326gat));
  OAI21_X1  g429(.A(G22gat), .B1(new_n591_), .B2(new_n547_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT42), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n547_), .A2(G22gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n606_), .B2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n333_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n315_), .A2(new_n254_), .A3(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(new_n590_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n638_), .A2(G29gat), .A3(new_n567_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n315_), .A2(new_n635_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n596_), .A2(KEYINPUT103), .A3(new_n597_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT103), .B1(new_n596_), .B2(new_n597_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n590_), .B2(KEYINPUT102), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n569_), .A2(new_n584_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n641_), .B1(new_n645_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n596_), .A2(new_n597_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n646_), .A2(KEYINPUT43), .A3(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT44), .B(new_n640_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT105), .ZN(new_n653_));
  INV_X1    g452(.A(new_n640_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n596_), .A2(KEYINPUT103), .A3(new_n597_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n511_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n549_), .B1(new_n661_), .B2(new_n558_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n567_), .B(new_n566_), .C1(new_n662_), .C2(new_n551_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n583_), .B1(new_n663_), .B2(new_n548_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n586_), .A2(new_n550_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(new_n547_), .A3(new_n588_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n664_), .A2(new_n666_), .A3(KEYINPUT102), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n659_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n651_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n654_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n671_), .A3(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n653_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT104), .B1(new_n670_), .B2(KEYINPUT44), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n664_), .B2(new_n666_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n648_), .A2(new_n677_), .A3(new_n658_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n651_), .B1(new_n678_), .B2(KEYINPUT43), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n675_), .B(new_n676_), .C1(new_n679_), .C2(new_n654_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n673_), .A2(new_n681_), .A3(new_n378_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G29gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G29gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n639_), .B1(new_n684_), .B2(new_n685_), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n673_), .A2(new_n681_), .A3(new_n560_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G36gat), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n638_), .A2(G36gat), .A3(new_n665_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n689_), .A2(KEYINPUT45), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(KEYINPUT45), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n688_), .A2(KEYINPUT46), .A3(new_n692_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n687_), .A2(G36gat), .B1(new_n691_), .B2(new_n690_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(G1329gat));
  NAND4_X1  g495(.A1(new_n673_), .A2(new_n681_), .A3(G43gat), .A4(new_n583_), .ZN(new_n697_));
  INV_X1    g496(.A(G43gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n638_), .B2(new_n584_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT47), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n697_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1330gat));
  AOI21_X1  g503(.A(G50gat), .B1(new_n637_), .B2(new_n566_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n673_), .A2(new_n681_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n566_), .A2(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(G1331gat));
  NOR3_X1   g507(.A1(new_n646_), .A2(new_n288_), .A3(new_n314_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n333_), .A2(new_n255_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n567_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n599_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT108), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n567_), .A2(G57gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n711_), .B2(new_n665_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n665_), .A2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n715_), .B2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n711_), .B2(new_n584_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n714_), .A2(new_n574_), .A3(new_n583_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n711_), .B2(new_n547_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT109), .Z(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT50), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT50), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n715_), .A2(G78gat), .A3(new_n547_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n288_), .A2(new_n635_), .A3(new_n314_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n679_), .B2(KEYINPUT111), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(KEYINPUT111), .B2(new_n679_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n567_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n709_), .A2(new_n255_), .A3(new_n333_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT110), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n738_), .A2(G85gat), .A3(new_n567_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g540(.A(G92gat), .B1(new_n735_), .B2(new_n665_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n665_), .A2(G92gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n738_), .B2(new_n743_), .ZN(G1337gat));
  OAI21_X1  g543(.A(G99gat), .B1(new_n735_), .B2(new_n584_), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n738_), .A2(new_n584_), .A3(new_n207_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g547(.A1(new_n738_), .A2(G106gat), .A3(new_n547_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n732_), .A2(new_n566_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n679_), .A2(KEYINPUT113), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT113), .B1(new_n679_), .B2(new_n751_), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n750_), .A2(new_n753_), .A3(new_n754_), .A4(G106gat), .ZN(new_n755_));
  INV_X1    g554(.A(G106gat), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n752_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n750_), .B1(new_n757_), .B2(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n749_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n749_), .C1(new_n755_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  AOI21_X1  g562(.A(new_n314_), .B1(KEYINPUT114), .B2(KEYINPUT54), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n288_), .A2(new_n635_), .A3(new_n650_), .A4(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n272_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n256_), .A2(new_n265_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n271_), .A2(new_n268_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(new_n267_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT115), .B(new_n274_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n267_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n769_), .A2(new_n774_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n283_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n283_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(KEYINPUT117), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n305_), .A2(new_n306_), .A3(new_n301_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n313_), .B1(new_n300_), .B2(new_n307_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n310_), .A2(new_n313_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n286_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n283_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n782_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n782_), .A2(KEYINPUT58), .A3(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n598_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n287_), .A2(new_n785_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT116), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n287_), .A2(new_n797_), .A3(new_n785_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n314_), .A2(new_n286_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n254_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT57), .B(new_n254_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n794_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n767_), .B1(new_n806_), .B2(new_n333_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n587_), .A2(new_n378_), .A3(new_n583_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n314_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n811_), .B1(KEYINPUT119), .B2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(KEYINPUT119), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(KEYINPUT119), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n807_), .A2(new_n810_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n815_), .A2(new_n314_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n819_), .B2(new_n812_), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n288_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n811_), .B(new_n822_), .C1(KEYINPUT60), .C2(new_n821_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT120), .ZN(new_n824_));
  INV_X1    g623(.A(new_n288_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n815_), .A2(new_n825_), .A3(new_n818_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n821_), .B2(new_n826_), .ZN(G1341gat));
  NAND4_X1  g626(.A1(new_n815_), .A2(G127gat), .A3(new_n635_), .A4(new_n818_), .ZN(new_n828_));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  INV_X1    g628(.A(new_n811_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n333_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n828_), .A2(KEYINPUT121), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT121), .B1(new_n828_), .B2(new_n831_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n811_), .A2(new_n835_), .A3(new_n255_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n815_), .A2(new_n598_), .A3(new_n818_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n835_), .ZN(G1343gat));
  NOR4_X1   g637(.A1(new_n560_), .A2(new_n583_), .A3(new_n567_), .A4(new_n547_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n807_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n314_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n825_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n635_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  AND3_X1   g647(.A1(new_n841_), .A2(G162gat), .A3(new_n658_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G162gat), .B1(new_n841_), .B2(new_n255_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n807_), .A2(new_n665_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n547_), .A3(new_n588_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n314_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n854_), .B(new_n855_), .C1(new_n859_), .C2(new_n429_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n429_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n861_));
  OAI221_X1 g660(.A(new_n861_), .B1(KEYINPUT123), .B2(KEYINPUT62), .C1(new_n857_), .C2(new_n858_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n862_), .A3(new_n863_), .ZN(G1348gat));
  NOR2_X1   g663(.A1(new_n857_), .A2(new_n288_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n428_), .A2(KEYINPUT124), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n428_), .A2(KEYINPUT124), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n865_), .B2(new_n867_), .ZN(G1349gat));
  NOR2_X1   g668(.A1(new_n857_), .A2(new_n333_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n410_), .A2(KEYINPUT125), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n411_), .A3(new_n413_), .A4(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT125), .A2(G183gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n870_), .B2(new_n873_), .ZN(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n857_), .B2(new_n650_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n255_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n857_), .B2(new_n876_), .ZN(G1351gat));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n568_), .A2(new_n583_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n856_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n878_), .B(new_n879_), .C1(new_n881_), .C2(new_n858_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n880_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n807_), .A2(new_n665_), .A3(new_n858_), .A4(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT127), .B1(new_n884_), .B2(KEYINPUT126), .ZN(new_n885_));
  AOI21_X1  g684(.A(G197gat), .B1(new_n884_), .B2(KEYINPUT126), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n882_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1352gat));
  AOI211_X1 g688(.A(new_n288_), .B(new_n881_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n881_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G204gat), .B1(new_n891_), .B2(new_n825_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1353gat));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  AND2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NOR4_X1   g694(.A1(new_n881_), .A2(new_n333_), .A3(new_n894_), .A4(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(new_n635_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n894_), .ZN(G1354gat));
  OR3_X1    g697(.A1(new_n881_), .A2(G218gat), .A3(new_n254_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G218gat), .B1(new_n881_), .B2(new_n650_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1355gat));
endmodule


