//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT67), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n212_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT6), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n211_), .A2(new_n213_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT10), .B(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n206_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n226_), .B(new_n227_), .C1(G85gat), .C2(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n215_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n217_), .A2(KEYINPUT8), .A3(new_n218_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n221_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n235_));
  XOR2_X1   g034(.A(G71gat), .B(G78gat), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n221_), .A2(new_n230_), .A3(new_n239_), .A4(new_n231_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n241_), .A2(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n203_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n241_), .A2(KEYINPUT12), .A3(new_n244_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT12), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n232_), .A2(new_n249_), .A3(new_n240_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n202_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G120gat), .B(G148gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT5), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G176gat), .B(G204gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n247_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(KEYINPUT13), .A3(new_n260_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT69), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G190gat), .B(G218gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT72), .ZN(new_n269_));
  XOR2_X1   g068(.A(G134gat), .B(G162gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G29gat), .B(G36gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT70), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G43gat), .B(G50gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n272_), .A2(KEYINPUT70), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(KEYINPUT70), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n281_), .A2(new_n221_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT34), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT35), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n280_), .B(KEYINPUT15), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n221_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n282_), .B(new_n287_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT15), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n280_), .B(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n293_), .B2(new_n232_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n285_), .A2(new_n286_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n290_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n232_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(new_n291_), .A3(new_n295_), .A4(new_n282_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n271_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT36), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT73), .B1(new_n297_), .B2(new_n299_), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT36), .B1(new_n305_), .B2(new_n271_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(new_n271_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT37), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT37), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G231gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n239_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G1gat), .ZN(new_n316_));
  INV_X1    g115(.A(G8gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT14), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G15gat), .B(G22gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G8gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT75), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n323_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n315_), .B(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G155gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G183gat), .B(G211gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT17), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n332_), .B(KEYINPUT17), .Z(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n327_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n313_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n326_), .A2(new_n280_), .ZN(new_n340_));
  AOI211_X1 g139(.A(new_n339_), .B(new_n340_), .C1(new_n293_), .C2(new_n326_), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n323_), .B(new_n325_), .Z(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n281_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n326_), .A2(new_n280_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT77), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n347_), .A3(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n341_), .B1(new_n349_), .B2(new_n339_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G141gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G169gat), .B(G197gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n350_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT82), .B1(new_n355_), .B2(KEYINPUT1), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(G155gat), .A4(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(G155gat), .B2(G162gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n355_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n365_), .A2(new_n366_), .B1(G141gat), .B2(G148gat), .ZN(new_n367_));
  INV_X1    g166(.A(G141gat), .ZN(new_n368_));
  INV_X1    g167(.A(G148gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(KEYINPUT3), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n374_), .A2(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT83), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n373_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n355_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n363_), .A2(new_n367_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n386_));
  INV_X1    g185(.A(G127gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(G134gat), .ZN(new_n388_));
  INV_X1    g187(.A(G134gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(G127gat), .ZN(new_n390_));
  INV_X1    g189(.A(G113gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(G120gat), .ZN(new_n392_));
  INV_X1    g191(.A(G120gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(G113gat), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n388_), .A2(new_n390_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G127gat), .B(G134gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n385_), .A2(new_n386_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n363_), .A2(new_n367_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n381_), .A2(new_n384_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT95), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(new_n398_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT80), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n401_), .A2(new_n402_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n400_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n406_), .A2(new_n407_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n384_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n372_), .A2(new_n370_), .B1(new_n379_), .B2(KEYINPUT83), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n378_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n356_), .A2(new_n359_), .B1(new_n361_), .B2(new_n355_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n366_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n376_), .B1(new_n422_), .B2(new_n364_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n417_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT95), .A3(new_n403_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n416_), .B1(new_n426_), .B2(new_n400_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n410_), .B1(new_n408_), .B2(new_n416_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n411_), .B(new_n415_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT33), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n409_), .A2(KEYINPUT4), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n428_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n435_), .A2(KEYINPUT97), .A3(new_n411_), .A4(new_n415_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n433_), .A3(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G8gat), .B(G36gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT19), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n447_));
  INV_X1    g246(.A(G176gat), .ZN(new_n448_));
  INV_X1    g247(.A(G169gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT22), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT22), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G169gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n448_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G169gat), .A2(G176gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G183gat), .A2(G190gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT23), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G183gat), .ZN(new_n461_));
  INV_X1    g260(.A(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT93), .ZN(new_n466_));
  AND3_X1   g265(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT93), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n463_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n456_), .A2(new_n457_), .A3(new_n466_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n461_), .A2(KEYINPUT25), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G183gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n462_), .A2(KEYINPUT26), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT26), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(G190gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n469_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT24), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n481_), .A2(G169gat), .A3(G176gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G169gat), .A2(G176gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n457_), .A2(KEYINPUT24), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT91), .B1(new_n480_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n485_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n469_), .A4(new_n479_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n472_), .A2(new_n487_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494_));
  INV_X1    g293(.A(G204gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(G197gat), .ZN(new_n496_));
  INV_X1    g295(.A(G197gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT21), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(G197gat), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n495_), .A2(G197gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n497_), .A2(G204gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT21), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G218gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G211gat), .ZN(new_n506_));
  INV_X1    g305(.A(G211gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G218gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(new_n504_), .A3(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n496_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n499_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n447_), .B1(new_n493_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n460_), .A2(new_n464_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n473_), .A2(new_n475_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G190gat), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G169gat), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n520_), .A2(new_n490_), .B1(new_n465_), .B2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n511_), .A2(KEYINPUT87), .A3(new_n514_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT87), .B1(new_n511_), .B2(new_n514_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n446_), .B1(new_n516_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n524_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n525_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n523_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n497_), .A2(G204gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n500_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n509_), .B1(KEYINPUT21), .B2(new_n533_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n534_), .A2(new_n501_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n472_), .A2(new_n535_), .A3(new_n487_), .A4(new_n492_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n445_), .A2(new_n447_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n531_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n443_), .B1(new_n527_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n471_), .A2(new_n466_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n451_), .A2(G169gat), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n449_), .A2(KEYINPUT22), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT92), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n450_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n544_));
  AOI21_X1  g343(.A(G176gat), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n457_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n540_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n487_), .A2(new_n492_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n515_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT20), .A3(new_n526_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n445_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n536_), .A2(new_n537_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n531_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n442_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n410_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n415_), .B1(new_n409_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n410_), .B1(new_n425_), .B2(KEYINPUT4), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n427_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n539_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n415_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n433_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n411_), .B(new_n561_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT96), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n435_), .A2(new_n564_), .A3(new_n411_), .A4(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n437_), .A2(new_n559_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n429_), .B1(new_n409_), .B2(KEYINPUT4), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n555_), .B1(new_n426_), .B2(new_n400_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n560_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n430_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n520_), .A2(new_n490_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n472_), .A2(new_n572_), .A3(new_n535_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n524_), .A2(new_n525_), .A3(new_n523_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n445_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n549_), .A2(KEYINPUT20), .A3(new_n446_), .A4(new_n526_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n442_), .A2(KEYINPUT32), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n550_), .A2(new_n445_), .B1(new_n552_), .B2(new_n531_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n571_), .B(new_n581_), .C1(new_n583_), .C2(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n567_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G78gat), .B(G106gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G228gat), .A2(G233gat), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT29), .B1(new_n420_), .B2(new_n424_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n535_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT88), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n587_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n528_), .A2(new_n588_), .A3(new_n529_), .A4(new_n587_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT90), .B(new_n586_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT84), .B1(new_n385_), .B2(new_n591_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT84), .A4(new_n591_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G22gat), .B(G50gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n401_), .A2(new_n402_), .A3(new_n591_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT84), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n598_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n600_), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n603_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n606_), .A2(new_n600_), .A3(new_n607_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n607_), .B1(new_n606_), .B2(new_n600_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n587_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n515_), .B1(new_n592_), .B2(KEYINPUT88), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n588_), .A2(new_n589_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n586_), .A2(KEYINPUT90), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n595_), .A3(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n597_), .A2(new_n609_), .A3(new_n613_), .A4(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n586_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n586_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n622_), .A3(new_n595_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(KEYINPUT89), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n613_), .A2(new_n609_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT89), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(new_n586_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n624_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n585_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n539_), .A2(new_n554_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT27), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n579_), .A2(new_n443_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n582_), .B2(new_n442_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n579_), .A2(KEYINPUT99), .A3(new_n443_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n570_), .A2(new_n430_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n629_), .A2(new_n634_), .A3(new_n640_), .A4(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT100), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n640_), .A2(new_n634_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n621_), .A2(new_n623_), .A3(KEYINPUT89), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n627_), .A3(new_n625_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n571_), .B1(new_n647_), .B2(new_n620_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n631_), .A2(new_n643_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G227gat), .A2(G233gat), .ZN(new_n652_));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(G71gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(G99gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT78), .B(G43gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n523_), .B(KEYINPUT30), .Z(new_n659_));
  INV_X1    g458(.A(KEYINPUT79), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n661_), .B2(new_n658_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n417_), .B(KEYINPUT31), .Z(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n666_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n650_), .A2(new_n651_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n644_), .A2(new_n630_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n669_), .A3(new_n571_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n651_), .B1(new_n650_), .B2(new_n669_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n354_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n267_), .B(new_n337_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n316_), .A3(new_n571_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT38), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n310_), .B(KEYINPUT104), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n669_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n630_), .A2(new_n585_), .B1(new_n642_), .B2(KEYINPUT100), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n649_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n672_), .B1(new_n687_), .B2(new_n651_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n650_), .A2(new_n669_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT101), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n684_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n263_), .A2(new_n264_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(KEYINPUT103), .A3(new_n354_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694_));
  INV_X1    g493(.A(new_n354_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n265_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n336_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n691_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G1gat), .B1(new_n700_), .B2(new_n641_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n680_), .A2(new_n681_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n682_), .A2(new_n701_), .A3(new_n702_), .ZN(G1324gat));
  INV_X1    g502(.A(new_n644_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n679_), .A2(new_n317_), .A3(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G8gat), .B1(new_n700_), .B2(new_n644_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT39), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n708_), .B(new_n709_), .Z(G1325gat));
  OAI21_X1  g509(.A(G15gat), .B1(new_n700_), .B2(new_n669_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT41), .Z(new_n712_));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n713_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n679_), .A2(new_n653_), .A3(new_n685_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT107), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT107), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n714_), .A2(new_n715_), .A3(new_n717_), .A4(new_n718_), .ZN(G1326gat));
  INV_X1    g518(.A(G22gat), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n629_), .B(KEYINPUT108), .Z(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n679_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G22gat), .B1(new_n700_), .B2(new_n721_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT42), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1327gat));
  NAND2_X1  g525(.A1(new_n310_), .A2(new_n698_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n265_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n731_), .A2(G29gat), .A3(new_n641_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n313_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n733_), .B(new_n734_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n313_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n697_), .A2(new_n336_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(KEYINPUT44), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT44), .B1(new_n738_), .B2(new_n739_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(new_n571_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n743_), .A2(KEYINPUT110), .A3(G29gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT110), .B1(new_n743_), .B2(G29gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n732_), .B1(new_n744_), .B2(new_n745_), .ZN(G1328gat));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n644_), .A2(G36gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n730_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(new_n730_), .B2(new_n750_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n740_), .A2(new_n741_), .A3(new_n644_), .ZN(new_n755_));
  INV_X1    g554(.A(G36gat), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n747_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n752_), .A2(new_n753_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(KEYINPUT46), .C1(new_n756_), .C2(new_n755_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1329gat));
  XOR2_X1   g560(.A(KEYINPUT112), .B(G43gat), .Z(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n731_), .B2(new_n669_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n742_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n685_), .A2(G43gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g567(.A(G50gat), .B1(new_n730_), .B2(new_n722_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n629_), .A2(G50gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n742_), .B2(new_n770_), .ZN(G1331gat));
  INV_X1    g570(.A(G57gat), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n337_), .A2(new_n692_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT113), .Z(new_n774_));
  AOI21_X1  g573(.A(new_n354_), .B1(new_n688_), .B2(new_n690_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n776_), .B2(new_n641_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n691_), .A2(new_n695_), .A3(new_n267_), .A4(new_n336_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n778_), .A2(new_n772_), .A3(new_n641_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(KEYINPUT114), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(KEYINPUT114), .B2(new_n779_), .ZN(G1332gat));
  OAI21_X1  g580(.A(G64gat), .B1(new_n778_), .B2(new_n644_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT48), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n644_), .A2(G64gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT115), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n776_), .B2(new_n785_), .ZN(G1333gat));
  OAI21_X1  g585(.A(G71gat), .B1(new_n778_), .B2(new_n669_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT49), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n669_), .A2(G71gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n776_), .B2(new_n789_), .ZN(G1334gat));
  OAI21_X1  g589(.A(G78gat), .B1(new_n778_), .B2(new_n721_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n721_), .A2(G78gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n776_), .B2(new_n794_), .ZN(G1335gat));
  NOR2_X1   g594(.A1(new_n266_), .A2(new_n727_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n775_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(G85gat), .B1(new_n798_), .B2(new_n571_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n265_), .A2(new_n695_), .A3(new_n698_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n733_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n737_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n800_), .B1(new_n803_), .B2(new_n735_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n571_), .A2(G85gat), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT117), .Z(new_n806_));
  AOI21_X1  g605(.A(new_n799_), .B1(new_n804_), .B2(new_n806_), .ZN(G1336gat));
  INV_X1    g606(.A(G92gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n797_), .B2(new_n644_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT118), .ZN(new_n810_));
  INV_X1    g609(.A(new_n804_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n811_), .A2(new_n808_), .A3(new_n644_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n811_), .B2(new_n669_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n798_), .A2(new_n685_), .A3(new_n224_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g616(.A(new_n800_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n738_), .A2(KEYINPUT119), .A3(new_n629_), .A4(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G106gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT119), .B1(new_n804_), .B2(new_n629_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n738_), .A2(new_n629_), .A3(new_n818_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(G106gat), .A4(new_n819_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n798_), .A2(new_n206_), .A3(new_n629_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  NOR3_X1   g633(.A1(new_n671_), .A2(new_n669_), .A3(new_n641_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n350_), .A2(new_n353_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n349_), .A2(new_n338_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n293_), .A2(new_n326_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n340_), .A2(new_n338_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n353_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n837_), .A2(new_n260_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n248_), .A2(new_n203_), .A3(new_n250_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n252_), .A2(KEYINPUT55), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n203_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n259_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n845_), .A2(KEYINPUT56), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n845_), .B2(new_n848_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n843_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n843_), .B(KEYINPUT58), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n309_), .A2(new_n853_), .A3(new_n312_), .A4(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n354_), .B(new_n260_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n261_), .A2(new_n837_), .A3(new_n842_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n859_), .B2(new_n308_), .ZN(new_n860_));
  AOI211_X1 g659(.A(KEYINPUT57), .B(new_n310_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n855_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT120), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n855_), .B(new_n864_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n698_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  AND4_X1   g666(.A1(new_n695_), .A2(new_n263_), .A3(new_n264_), .A4(new_n336_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n313_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n313_), .B2(new_n868_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n836_), .B1(new_n866_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n391_), .A3(new_n354_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n336_), .B1(new_n862_), .B2(KEYINPUT120), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n875_), .B2(new_n865_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n876_), .B2(new_n836_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n862_), .A2(new_n698_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n872_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n835_), .B2(KEYINPUT121), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(KEYINPUT121), .B2(new_n835_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n877_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n354_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n874_), .B1(new_n886_), .B2(new_n391_), .ZN(G1340gat));
  OAI211_X1 g686(.A(new_n883_), .B(new_n267_), .C1(new_n873_), .C2(new_n880_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n692_), .A2(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n873_), .B1(KEYINPUT60), .B2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n877_), .A2(KEYINPUT122), .A3(new_n267_), .A4(new_n883_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n890_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  OAI22_X1  g693(.A1(new_n894_), .A2(new_n393_), .B1(KEYINPUT60), .B2(new_n892_), .ZN(G1341gat));
  NAND3_X1  g694(.A1(new_n873_), .A2(new_n387_), .A3(new_n336_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n884_), .A2(new_n336_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n387_), .ZN(G1342gat));
  AOI21_X1  g698(.A(G134gat), .B1(new_n873_), .B2(new_n684_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n900_), .A2(KEYINPUT123), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(KEYINPUT123), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n313_), .A2(new_n389_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n901_), .A2(new_n902_), .B1(new_n884_), .B2(new_n903_), .ZN(G1343gat));
  NAND2_X1  g703(.A1(new_n629_), .A2(new_n571_), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n876_), .A2(new_n685_), .A3(new_n704_), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n354_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n267_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n336_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  INV_X1    g712(.A(G162gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n906_), .B2(new_n733_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n683_), .A2(G162gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n906_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(KEYINPUT124), .A3(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  INV_X1    g719(.A(new_n918_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n915_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n919_), .A2(new_n922_), .ZN(G1347gat));
  AOI21_X1  g722(.A(new_n722_), .B1(new_n872_), .B2(new_n878_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n704_), .A2(new_n641_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n669_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n354_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(G169gat), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n928_), .B(new_n354_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n930_), .B1(new_n929_), .B2(G169gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1348gat));
  AOI21_X1  g734(.A(G176gat), .B1(new_n928_), .B2(new_n265_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n876_), .A2(new_n629_), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n266_), .A2(new_n448_), .A3(new_n669_), .A4(new_n925_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n925_), .A2(new_n669_), .A3(new_n698_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G183gat), .B1(new_n937_), .B2(new_n940_), .ZN(new_n941_));
  NOR4_X1   g740(.A1(new_n925_), .A2(new_n518_), .A3(new_n669_), .A4(new_n698_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n924_), .B2(new_n942_), .ZN(G1350gat));
  NAND2_X1  g742(.A1(new_n928_), .A2(new_n733_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(new_n945_), .A3(G190gat), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n944_), .B2(G190gat), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n684_), .A2(new_n519_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT126), .ZN(new_n950_));
  OAI22_X1  g749(.A1(new_n947_), .A2(new_n948_), .B1(new_n927_), .B2(new_n950_), .ZN(G1351gat));
  NOR2_X1   g750(.A1(new_n876_), .A2(new_n685_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n952_), .A2(new_n704_), .A3(new_n641_), .A4(new_n629_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n695_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(new_n497_), .ZN(G1352gat));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n266_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n956_), .B1(KEYINPUT127), .B2(new_n495_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(KEYINPUT127), .B(G204gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n956_), .B2(new_n958_), .ZN(G1353gat));
  NOR2_X1   g758(.A1(new_n953_), .A2(new_n698_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  AND2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n960_), .B1(new_n961_), .B2(new_n962_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(new_n960_), .B2(new_n961_), .ZN(G1354gat));
  OAI21_X1  g763(.A(G218gat), .B1(new_n953_), .B2(new_n313_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n684_), .A2(new_n505_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n953_), .B2(new_n966_), .ZN(G1355gat));
endmodule


