//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT80), .Z(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT1), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n209_), .B(new_n210_), .C1(new_n212_), .C2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n211_), .B(KEYINPUT80), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT3), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n210_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT81), .B(KEYINPUT2), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n210_), .B1(KEYINPUT81), .B2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n216_), .B(new_n213_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n215_), .A2(new_n226_), .A3(KEYINPUT82), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT82), .B1(new_n215_), .B2(new_n226_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n206_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n215_), .A2(new_n226_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(new_n206_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n230_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n231_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(new_n227_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n232_), .B1(new_n242_), .B2(new_n206_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n239_), .B1(new_n243_), .B2(new_n238_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n237_), .B1(new_n244_), .B2(new_n236_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  OAI21_X1  g048(.A(new_n202_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n238_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT4), .B1(new_n242_), .B2(new_n206_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n236_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n237_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n249_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT94), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n254_), .A3(new_n249_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT23), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(G183gat), .B2(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT76), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT22), .B(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n263_), .B(new_n264_), .C1(new_n265_), .C2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n265_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G190gat), .ZN(new_n273_));
  INV_X1    g072(.A(G183gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT25), .B1(new_n274_), .B2(KEYINPUT74), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n274_), .A2(KEYINPUT25), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n275_), .C1(new_n276_), .C2(KEYINPUT74), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT75), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n262_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n286_), .A3(new_n280_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n272_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G197gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(G204gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT84), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT84), .ZN(new_n293_));
  INV_X1    g092(.A(G204gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(G197gat), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n292_), .B(KEYINPUT21), .C1(new_n291_), .C2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G211gat), .B(G218gat), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n290_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT85), .B1(new_n290_), .B2(G204gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(new_n291_), .B2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n296_), .B(new_n298_), .C1(new_n301_), .C2(KEYINPUT21), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT21), .A3(new_n297_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n260_), .B1(new_n289_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n264_), .B(KEYINPUT89), .Z(new_n307_));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n266_), .B(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n263_), .B(new_n307_), .C1(new_n309_), .C2(G176gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n273_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT25), .B(G183gat), .Z(new_n312_));
  OAI211_X1 g111(.A(new_n285_), .B(new_n280_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT88), .ZN(new_n317_));
  XOR2_X1   g116(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n272_), .A2(new_n288_), .A3(new_n306_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n310_), .A2(new_n313_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n260_), .B1(new_n322_), .B2(new_n304_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n320_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n324_), .A2(new_n319_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n288_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n269_), .A2(new_n271_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n304_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n319_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n337_), .A2(KEYINPUT20), .A3(new_n338_), .A4(new_n314_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n340_), .A2(new_n332_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n259_), .A2(new_n333_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n330_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n334_), .A2(new_n331_), .A3(new_n339_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n334_), .A2(new_n339_), .A3(KEYINPUT92), .A4(new_n331_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n234_), .A2(new_n235_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n244_), .B2(new_n235_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n346_), .A2(new_n347_), .B1(new_n256_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n258_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT33), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n258_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n342_), .A2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n205_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT79), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT77), .ZN(new_n364_));
  XOR2_X1   g163(.A(G15gat), .B(G43gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n361_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G71gat), .B(G99gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n289_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n361_), .A2(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n361_), .A2(new_n366_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n228_), .A2(new_n229_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT28), .B1(new_n242_), .B2(KEYINPUT29), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(G228gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(G228gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(new_n304_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n231_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n396_));
  OAI21_X1  g195(.A(new_n304_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n392_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n394_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n386_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n405_), .A2(new_n385_), .A3(new_n383_), .A4(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n357_), .A2(new_n375_), .A3(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n404_), .A2(new_n375_), .A3(new_n406_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n375_), .B1(new_n406_), .B2(new_n404_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n259_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n346_), .A2(new_n414_), .A3(new_n347_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n325_), .A2(new_n330_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT27), .A3(new_n345_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n408_), .B1(new_n411_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT68), .ZN(new_n420_));
  INV_X1    g219(.A(G57gat), .ZN(new_n421_));
  INV_X1    g220(.A(G64gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G57gat), .A2(G64gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT11), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G78gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n423_), .A2(new_n429_), .A3(new_n424_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n427_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G85gat), .B(G92gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT7), .ZN(new_n434_));
  INV_X1    g233(.A(G99gat), .ZN(new_n435_));
  INV_X1    g234(.A(G106gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n433_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT67), .B1(new_n441_), .B2(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  NAND3_X1  g249(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n439_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n433_), .A2(KEYINPUT8), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n444_), .A2(new_n445_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G85gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT66), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G85gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n458_), .A2(new_n460_), .A3(G92gat), .A4(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n457_), .A2(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(G92gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n446_), .A2(new_n452_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT10), .B(G99gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n471_), .B2(G106gat), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n435_), .A2(KEYINPUT10), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n435_), .A2(KEYINPUT10), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT64), .B(new_n436_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n469_), .A3(new_n472_), .A4(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n432_), .B1(new_n456_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n420_), .B(KEYINPUT12), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT67), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n450_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n440_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n454_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n433_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n449_), .A2(new_n451_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n484_), .B1(new_n439_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT8), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n464_), .A2(new_n467_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n472_), .A2(new_n475_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n483_), .A2(new_n487_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n432_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n479_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n420_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT12), .B1(new_n477_), .B2(new_n420_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n428_), .A2(new_n431_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n462_), .A2(new_n463_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n480_), .A2(new_n481_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n489_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n482_), .A2(new_n454_), .B1(new_n486_), .B2(KEYINPUT8), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n492_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n494_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT5), .B(G176gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G204gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n498_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n498_), .B2(new_n507_), .ZN(new_n515_));
  AND2_X1   g314(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n516_));
  OR3_X1    g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n518_));
  OAI22_X1  g317(.A1(new_n514_), .A2(new_n515_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G15gat), .B(G22gat), .Z(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT73), .B(G1gat), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G8gat), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n523_), .B2(KEYINPUT14), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G29gat), .B(G36gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G43gat), .B(G50gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n524_), .A2(new_n525_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n525_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n529_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n540_));
  NOR2_X1   g339(.A1(new_n529_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n539_), .B1(new_n542_), .B2(new_n538_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n539_), .B(new_n548_), .C1(new_n542_), .C2(new_n538_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n520_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n419_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n526_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n432_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G127gat), .B(G155gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G211gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT16), .B(G183gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT17), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(KEYINPUT17), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n556_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n562_), .B2(new_n556_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n540_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n530_), .B1(new_n491_), .B2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n540_), .B(new_n529_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT72), .ZN(new_n574_));
  INV_X1    g373(.A(G232gat), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(new_n387_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n573_), .A2(KEYINPUT72), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n579_), .A3(KEYINPUT34), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT34), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n573_), .B2(KEYINPUT72), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n583_));
  AOI211_X1 g382(.A(new_n583_), .B(new_n576_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT35), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n573_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n580_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT35), .B1(new_n580_), .B2(new_n585_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n566_), .B(new_n569_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n580_), .A2(new_n585_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n586_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n569_), .A2(new_n566_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n569_), .A2(new_n566_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n580_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n590_), .A2(new_n596_), .A3(KEYINPUT37), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n553_), .A2(new_n565_), .A3(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT96), .Z(new_n604_));
  INV_X1    g403(.A(new_n522_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n259_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT97), .Z(new_n609_));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n597_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n590_), .A2(new_n596_), .A3(KEYINPUT98), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n565_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n553_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n259_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n606_), .A2(new_n607_), .B1(G1gat), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n609_), .A2(new_n618_), .ZN(G1324gat));
  AND2_X1   g418(.A1(new_n417_), .A2(new_n415_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G8gat), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT39), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n623_), .B(KEYINPUT99), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(G8gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n604_), .A2(new_n630_), .A3(new_n621_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(G1325gat));
  INV_X1    g433(.A(G15gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n375_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n604_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n635_), .B1(new_n616_), .B2(new_n636_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1326gat));
  INV_X1    g439(.A(G22gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n407_), .B(KEYINPUT101), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n616_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n604_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1327gat));
  AND3_X1   g445(.A1(new_n590_), .A2(new_n596_), .A3(KEYINPUT98), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT98), .B1(new_n590_), .B2(new_n596_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n565_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n553_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT104), .Z(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n259_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  INV_X1    g453(.A(new_n407_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n636_), .B(new_n655_), .C1(new_n342_), .C2(new_n356_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n418_), .A2(new_n411_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n601_), .B(new_n654_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n656_), .A2(new_n657_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n661_), .B2(new_n602_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n419_), .A2(KEYINPUT102), .A3(new_n654_), .A4(new_n601_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n552_), .A3(new_n614_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n664_), .A2(KEYINPUT44), .A3(new_n552_), .A4(new_n614_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n669_), .A2(KEYINPUT103), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT103), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n259_), .A2(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n653_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n652_), .A2(new_n676_), .A3(new_n621_), .ZN(new_n677_));
  XOR2_X1   g476(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n678_));
  XOR2_X1   g477(.A(new_n677_), .B(new_n678_), .Z(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n672_), .B2(new_n621_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n680_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n677_), .B(new_n678_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1329gat));
  NAND2_X1  g484(.A1(new_n652_), .A2(new_n636_), .ZN(new_n686_));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n375_), .A2(new_n687_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n672_), .B2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n669_), .A2(KEYINPUT103), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n669_), .A2(KEYINPUT103), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n667_), .B(new_n690_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(KEYINPUT106), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n688_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT47), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(new_n688_), .C1(new_n691_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1330gat));
  AOI21_X1  g499(.A(G50gat), .B1(new_n652_), .B2(new_n642_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n672_), .A2(G50gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n703_), .B2(new_n655_), .ZN(G1331gat));
  INV_X1    g503(.A(new_n520_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n550_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n419_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n601_), .A2(new_n614_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n421_), .B1(new_n709_), .B2(new_n412_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n615_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n259_), .A2(G57gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT107), .ZN(G1332gat));
  OAI21_X1  g513(.A(G64gat), .B1(new_n711_), .B2(new_n620_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT48), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n621_), .A2(new_n422_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n709_), .B2(new_n717_), .ZN(G1333gat));
  OAI21_X1  g517(.A(G71gat), .B1(new_n711_), .B2(new_n375_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT49), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n375_), .A2(G71gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n709_), .B2(new_n721_), .ZN(G1334gat));
  INV_X1    g521(.A(new_n642_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G78gat), .B1(new_n711_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT50), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n723_), .A2(G78gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n709_), .B2(new_n726_), .ZN(G1335gat));
  NAND2_X1  g526(.A1(new_n707_), .A2(new_n650_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n259_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n664_), .A2(new_n614_), .A3(new_n706_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n259_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(G1336gat));
  AOI21_X1  g532(.A(G92gat), .B1(new_n729_), .B2(new_n621_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n731_), .A2(new_n621_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G92gat), .ZN(G1337gat));
  OR3_X1    g535(.A1(new_n728_), .A2(new_n471_), .A3(new_n375_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n731_), .A2(new_n636_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n435_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n740_));
  OR2_X1    g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n741_), .A2(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(KEYINPUT51), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(KEYINPUT109), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n729_), .A2(new_n436_), .A3(new_n655_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n731_), .A2(new_n655_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G106gat), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT52), .B(new_n436_), .C1(new_n731_), .C2(new_n655_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g551(.A1(new_n621_), .A2(new_n412_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n410_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n536_), .A2(new_n537_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n546_), .C1(new_n542_), .C2(new_n537_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n549_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n758_), .B(KEYINPUT111), .C1(new_n514_), .C2(new_n515_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT68), .B1(new_n504_), .B2(KEYINPUT69), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT12), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n504_), .B2(KEYINPUT68), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n492_), .B(new_n479_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n765_), .B1(new_n769_), .B2(new_n506_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n506_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n769_), .A2(new_n765_), .A3(new_n506_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n511_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n764_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n494_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n498_), .B1(new_n777_), .B2(new_n765_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n773_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n512_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT56), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n551_), .B1(new_n776_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n764_), .A3(KEYINPUT56), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n513_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n763_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT112), .B1(new_n785_), .B2(new_n613_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  INV_X1    g586(.A(new_n763_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT110), .B1(new_n780_), .B2(KEYINPUT56), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n775_), .B(new_n512_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n550_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n783_), .A2(new_n513_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n649_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n786_), .A2(new_n787_), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT57), .A3(new_n649_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n774_), .A2(new_n775_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n781_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n514_), .B1(new_n790_), .B2(KEYINPUT113), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n758_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT114), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT58), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(KEYINPUT114), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n601_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n796_), .A2(new_n797_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n796_), .A2(new_n807_), .A3(KEYINPUT115), .A4(new_n797_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n614_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n708_), .A2(new_n551_), .A3(new_n705_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT54), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n755_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815_), .B2(new_n550_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n796_), .A2(new_n817_), .A3(new_n807_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n797_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n796_), .B2(new_n807_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n614_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n814_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n755_), .A2(KEYINPUT59), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n815_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n551_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n816_), .B1(new_n827_), .B2(G113gat), .ZN(G1340gat));
  XNOR2_X1  g627(.A(KEYINPUT118), .B(G120gat), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n705_), .B2(new_n829_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n815_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n832_), .B2(new_n830_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n826_), .A2(new_n832_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n520_), .ZN(G1341gat));
  AOI21_X1  g634(.A(G127gat), .B1(new_n815_), .B2(new_n565_), .ZN(new_n836_));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n826_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n565_), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n602_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n824_), .B(new_n841_), .C1(new_n825_), .C2(new_n815_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n649_), .B(new_n755_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT119), .B1(new_n843_), .B2(G134gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n815_), .A2(new_n613_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n840_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n844_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n842_), .A2(new_n844_), .A3(new_n847_), .A4(KEYINPUT120), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1343gat));
  NAND2_X1  g651(.A1(new_n812_), .A2(new_n814_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n409_), .A3(new_n753_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n551_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n207_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n705_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT121), .B(G148gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1345gat));
  NOR2_X1   g658(.A1(new_n854_), .A2(new_n614_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT61), .B(G155gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n854_), .A2(new_n649_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(G162gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n601_), .A2(G162gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT122), .Z(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n854_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n863_), .B1(new_n865_), .B2(new_n869_), .ZN(new_n870_));
  OAI221_X1 g669(.A(KEYINPUT123), .B1(new_n854_), .B2(new_n868_), .C1(new_n864_), .C2(G162gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1347gat));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n620_), .A2(new_n259_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n636_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n642_), .A2(new_n551_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n822_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(G169gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n873_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n875_), .B1(new_n821_), .B2(new_n814_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n877_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(KEYINPUT62), .A3(new_n883_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n882_), .A2(new_n309_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n873_), .B(new_n886_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .ZN(G1348gat));
  AND2_X1   g687(.A1(new_n881_), .A2(new_n723_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G176gat), .B1(new_n889_), .B2(new_n520_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n655_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n875_), .A2(new_n705_), .A3(new_n267_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1349gat));
  NAND4_X1  g692(.A1(new_n881_), .A2(new_n312_), .A3(new_n565_), .A4(new_n723_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n895_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n875_), .A2(new_n614_), .ZN(new_n898_));
  AOI21_X1  g697(.A(G183gat), .B1(new_n891_), .B2(new_n898_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n896_), .A2(new_n897_), .A3(new_n899_), .ZN(G1350gat));
  NAND2_X1  g699(.A1(new_n889_), .A2(new_n601_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G190gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n889_), .A2(new_n273_), .A3(new_n613_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1351gat));
  NAND3_X1  g703(.A1(new_n853_), .A2(new_n409_), .A3(new_n874_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT126), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n853_), .A2(new_n907_), .A3(new_n409_), .A4(new_n874_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G197gat), .B1(new_n909_), .B2(new_n550_), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n290_), .B(new_n551_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1352gat));
  AOI21_X1  g711(.A(G204gat), .B1(new_n909_), .B2(new_n520_), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n294_), .B(new_n705_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1353gat));
  OR2_X1    g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n909_), .B2(new_n565_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  AOI211_X1 g717(.A(new_n614_), .B(new_n918_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1354gat));
  XOR2_X1   g719(.A(KEYINPUT127), .B(G218gat), .Z(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n909_), .B2(new_n613_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n602_), .B(new_n923_), .C1(new_n906_), .C2(new_n908_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1355gat));
endmodule


