//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n207_), .A2(KEYINPUT2), .B1(new_n210_), .B2(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT89), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n206_), .B(new_n212_), .ZN(new_n213_));
  OAI221_X1 g012(.A(new_n211_), .B1(KEYINPUT3), .B2(new_n210_), .C1(new_n213_), .C2(KEYINPUT2), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT90), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n217_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n215_), .B(KEYINPUT1), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n210_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n213_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT99), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n205_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n223_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G225gat), .A2(G233gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n226_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n204_), .A2(KEYINPUT4), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n229_), .A2(KEYINPUT4), .B1(new_n222_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n228_), .B1(new_n231_), .B2(new_n227_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G1gat), .B(G29gat), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G57gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT33), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G183gat), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT23), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT85), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT85), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT23), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G183gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n242_), .A2(KEYINPUT25), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .A4(new_n257_), .ZN(new_n258_));
  OR3_X1    g057(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT84), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n250_), .A2(new_n258_), .A3(new_n259_), .A4(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n249_), .A2(new_n244_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(G183gat), .B2(G190gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(G176gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(new_n261_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G197gat), .B(G204gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n274_), .A2(new_n275_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n273_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n248_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n271_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n263_), .A2(new_n260_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n255_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n266_), .A2(new_n259_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n284_), .B1(new_n292_), .B2(new_n282_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n283_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G64gat), .B(G92gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G8gat), .B(G36gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n296_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT20), .B(new_n304_), .C1(new_n292_), .C2(new_n282_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT96), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n273_), .A2(new_n307_), .A3(new_n282_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(new_n273_), .B2(new_n282_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n306_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n297_), .A2(new_n303_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n273_), .A2(new_n282_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT96), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n305_), .B1(new_n314_), .B2(new_n308_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n304_), .B1(new_n283_), .B2(new_n293_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n302_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n317_), .A3(KEYINPUT98), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT98), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n297_), .A2(new_n311_), .A3(new_n319_), .A4(new_n303_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n231_), .A2(new_n227_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n237_), .C1(new_n227_), .C2(new_n226_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n232_), .A2(KEYINPUT33), .A3(new_n238_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n241_), .A2(new_n321_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n294_), .A2(new_n296_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n282_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n280_), .A2(KEYINPUT92), .A3(new_n281_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI221_X1 g129(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n292_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n331_), .B2(new_n296_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n297_), .A2(new_n311_), .A3(new_n333_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n232_), .A2(new_n238_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n232_), .A2(new_n238_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n334_), .B(new_n335_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n325_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT30), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n273_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n342_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT86), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n344_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n345_), .B1(new_n344_), .B2(new_n351_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n204_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n205_), .A3(new_n352_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n343_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n357_), .A3(new_n343_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(KEYINPUT88), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT88), .ZN(new_n362_));
  INV_X1    g161(.A(new_n360_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT94), .ZN(new_n366_));
  AOI22_X1  g165(.A1(KEYINPUT29), .A2(new_n222_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n370_), .A2(new_n368_), .A3(new_n282_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n373_), .B(KEYINPUT93), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n370_), .A2(new_n368_), .A3(new_n282_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(KEYINPUT94), .C1(new_n368_), .C2(new_n367_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT95), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n369_), .A2(new_n371_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n374_), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n222_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT28), .B(G22gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(G50gat), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n384_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n372_), .A2(KEYINPUT95), .A3(new_n375_), .A4(new_n377_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n380_), .A2(new_n382_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(KEYINPUT91), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n382_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n381_), .A2(new_n374_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n392_), .B(new_n394_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n391_), .A2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n339_), .A2(new_n365_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT27), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n318_), .A2(new_n400_), .A3(new_n320_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT27), .B(new_n312_), .C1(new_n332_), .C2(new_n303_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n398_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT101), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n359_), .A2(new_n360_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT101), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n398_), .B(new_n409_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n398_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n365_), .A2(new_n412_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n337_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n239_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n399_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G176gat), .B(G204gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G120gat), .B(G148gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  XOR2_X1   g223(.A(G85gat), .B(G92gat), .Z(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT10), .B(G99gat), .Z(new_n426_));
  INV_X1    g225(.A(G106gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(KEYINPUT9), .A2(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT64), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT6), .ZN(new_n432_));
  AND2_X1   g231(.A1(G99gat), .A2(G106gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n428_), .B(new_n436_), .C1(KEYINPUT9), .C2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT66), .B1(new_n434_), .B2(new_n435_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n433_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n431_), .A2(KEYINPUT6), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n429_), .A2(KEYINPUT64), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT7), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n439_), .B1(new_n450_), .B2(new_n425_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n446_), .A3(new_n444_), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n453_));
  AND3_X1   g252(.A1(new_n452_), .A2(new_n425_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n438_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(KEYINPUT68), .B(new_n438_), .C1(new_n451_), .C2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G64gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(KEYINPUT11), .ZN(new_n462_));
  XOR2_X1   g261(.A(G71gat), .B(G78gat), .Z(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n462_), .A2(new_n463_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT12), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n459_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G230gat), .A2(G233gat), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n438_), .B(new_n466_), .C1(new_n451_), .C2(new_n454_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT12), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n455_), .A2(new_n467_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(new_n472_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n471_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n478_), .B(new_n479_), .C1(new_n477_), .C2(new_n472_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n424_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n476_), .A2(new_n480_), .A3(new_n424_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT71), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n483_), .A2(KEYINPUT70), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n483_), .B2(KEYINPUT70), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(KEYINPUT70), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT71), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(KEYINPUT70), .A3(new_n484_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n481_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n487_), .A2(new_n491_), .B1(new_n492_), .B2(KEYINPUT13), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(KEYINPUT13), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT13), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n487_), .A2(new_n491_), .A3(KEYINPUT72), .A4(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G1gat), .B(G8gat), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT76), .B(G22gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(G15gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n504_));
  INV_X1    g303(.A(G1gat), .ZN(new_n505_));
  INV_X1    g304(.A(G8gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n503_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n501_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT77), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n503_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n500_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n510_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT79), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n510_), .A2(new_n514_), .A3(KEYINPUT79), .A4(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n514_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n517_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n526_), .A2(KEYINPUT80), .A3(G229gat), .A4(G233gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT80), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n520_), .A2(new_n521_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(KEYINPUT81), .ZN(new_n532_));
  INV_X1    g331(.A(new_n523_), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n517_), .B(KEYINPUT15), .Z(new_n534_));
  OAI211_X1 g333(.A(new_n522_), .B(new_n532_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n527_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n527_), .A2(new_n531_), .A3(new_n535_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n499_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n534_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n517_), .B(new_n438_), .C1(new_n451_), .C2(new_n454_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT73), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n548_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n546_), .A2(new_n459_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G232gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT34), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n554_), .A2(new_n555_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n551_), .A2(KEYINPUT35), .A3(new_n553_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(G162gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT74), .B(G134gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  AOI22_X1  g365(.A1(new_n560_), .A2(new_n561_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(new_n562_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n560_), .A2(new_n569_), .A3(new_n561_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n570_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n567_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n523_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n466_), .B(KEYINPUT78), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n578_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583_));
  INV_X1    g382(.A(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT16), .B(G183gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n582_), .B1(KEYINPUT17), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n587_), .B(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n591_), .B2(new_n582_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n576_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n419_), .A2(new_n545_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n505_), .A3(new_n416_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n574_), .A2(new_n567_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT102), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n419_), .A2(new_n545_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n417_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(G1324gat));
  NOR2_X1   g402(.A1(new_n404_), .A2(new_n405_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G8gat), .B1(new_n601_), .B2(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT103), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(KEYINPUT103), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(KEYINPUT104), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n595_), .A2(new_n506_), .A3(new_n604_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(KEYINPUT104), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n607_), .A2(new_n608_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n611_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n611_), .A2(KEYINPUT40), .A3(new_n612_), .A4(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n601_), .B2(new_n365_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT41), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n594_), .A2(G15gat), .A3(new_n365_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1326gat));
  OAI21_X1  g423(.A(G22gat), .B1(new_n601_), .B2(new_n398_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT42), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n398_), .A2(G22gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n594_), .B2(new_n627_), .ZN(G1327gat));
  NOR2_X1   g427(.A1(new_n418_), .A2(new_n598_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n545_), .A3(new_n592_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n630_), .A2(G29gat), .A3(new_n417_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n545_), .A2(new_n592_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n576_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT43), .B1(new_n418_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n416_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n635_), .B(new_n576_), .C1(new_n636_), .C2(new_n399_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n632_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT44), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n417_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n634_), .A2(new_n637_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n632_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT105), .A3(G29gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT105), .B1(new_n644_), .B2(G29gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n631_), .B1(new_n645_), .B2(new_n646_), .ZN(G1328gat));
  NOR3_X1   g446(.A1(new_n630_), .A2(G36gat), .A3(new_n605_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT45), .Z(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n605_), .B1(new_n638_), .B2(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n652_), .B2(G36gat), .ZN(new_n653_));
  INV_X1    g452(.A(G36gat), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT106), .B(new_n654_), .C1(new_n643_), .C2(new_n651_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n649_), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI221_X1 g457(.A(new_n649_), .B1(KEYINPUT107), .B2(KEYINPUT46), .C1(new_n653_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1329gat));
  NAND3_X1  g459(.A1(new_n643_), .A2(G43gat), .A3(new_n408_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n630_), .A2(new_n365_), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n661_), .A2(new_n639_), .B1(G43gat), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g463(.A1(new_n643_), .A2(new_n412_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G50gat), .B1(new_n665_), .B2(new_n639_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n398_), .A2(G50gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT108), .Z(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n630_), .B2(new_n668_), .ZN(G1331gat));
  NAND2_X1  g468(.A1(new_n499_), .A2(new_n544_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n418_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n600_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n417_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n593_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT109), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(KEYINPUT109), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n677_), .A2(KEYINPUT110), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT110), .B1(new_n677_), .B2(new_n678_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n416_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n674_), .B1(new_n681_), .B2(new_n673_), .ZN(G1332gat));
  NOR2_X1   g481(.A1(new_n677_), .A2(new_n678_), .ZN(new_n683_));
  INV_X1    g482(.A(G64gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n604_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G64gat), .B1(new_n672_), .B2(new_n605_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1333gat));
  OAI21_X1  g488(.A(G71gat), .B1(new_n672_), .B2(new_n365_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT49), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n365_), .A2(G71gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT112), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n683_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1334gat));
  INV_X1    g494(.A(G78gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n683_), .A2(new_n696_), .A3(new_n412_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G78gat), .B1(new_n672_), .B2(new_n398_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT50), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1335gat));
  INV_X1    g499(.A(new_n592_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n670_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n629_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n416_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n634_), .A2(new_n637_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n702_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n417_), .A2(new_n234_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(G1336gat));
  AOI21_X1  g508(.A(G92gat), .B1(new_n704_), .B2(new_n604_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n604_), .A2(G92gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n707_), .B2(new_n711_), .ZN(G1337gat));
  AND3_X1   g511(.A1(new_n704_), .A2(new_n426_), .A3(new_n408_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n365_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n707_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n715_), .B2(G99gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n706_), .A2(new_n412_), .A3(new_n702_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(new_n427_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(KEYINPUT52), .A3(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n704_), .A2(new_n427_), .A3(new_n412_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n718_), .B(new_n725_), .C1(new_n720_), .C2(new_n427_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT53), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT53), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n723_), .A2(new_n729_), .A3(new_n724_), .A4(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1339gat));
  INV_X1    g530(.A(new_n424_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n473_), .A2(new_n474_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n468_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n479_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n479_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(KEYINPUT55), .B2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n470_), .A2(KEYINPUT55), .A3(new_n471_), .A4(new_n475_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n732_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT56), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n526_), .A2(new_n532_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n532_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n522_), .B(new_n743_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(new_n539_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n742_), .A2(KEYINPUT114), .A3(new_n744_), .A4(new_n539_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n542_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n471_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n476_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n738_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n732_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n741_), .A2(new_n749_), .A3(new_n483_), .A4(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT58), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n754_), .B1(new_n753_), .B2(new_n732_), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT56), .B(new_n424_), .C1(new_n752_), .C2(new_n738_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT58), .A3(new_n483_), .A4(new_n749_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(new_n762_), .A3(new_n576_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT115), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n741_), .A2(new_n543_), .A3(new_n483_), .A4(new_n755_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n487_), .A2(new_n491_), .A3(new_n749_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT57), .A3(new_n598_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n598_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n758_), .A2(new_n762_), .A3(new_n576_), .A4(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n764_), .A2(new_n768_), .A3(new_n771_), .A4(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n592_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n593_), .A2(new_n544_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT54), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n411_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n777_), .A3(KEYINPUT116), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n780_), .A2(new_n416_), .A3(new_n781_), .A4(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G113gat), .B1(new_n784_), .B2(new_n543_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(KEYINPUT59), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n771_), .A2(new_n768_), .A3(new_n763_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n592_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n777_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n417_), .A2(KEYINPUT59), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n781_), .A3(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT118), .Z(new_n794_));
  NAND3_X1  g593(.A1(new_n783_), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n788_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n543_), .A2(G113gat), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT119), .Z(new_n798_));
  AOI21_X1  g597(.A(new_n785_), .B1(new_n796_), .B2(new_n798_), .ZN(G1340gat));
  NAND4_X1  g598(.A1(new_n788_), .A2(new_n794_), .A3(new_n499_), .A4(new_n795_), .ZN(new_n800_));
  INV_X1    g599(.A(G120gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT60), .B1(new_n499_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n783_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G120gat), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n803_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(KEYINPUT60), .B2(new_n805_), .ZN(G1341gat));
  AOI21_X1  g605(.A(G127gat), .B1(new_n784_), .B2(new_n701_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n701_), .A2(G127gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n796_), .B2(new_n808_), .ZN(G1342gat));
  NAND2_X1  g608(.A1(new_n576_), .A2(G134gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT120), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n788_), .A2(new_n794_), .A3(new_n795_), .A4(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  INV_X1    g612(.A(new_n599_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n783_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT121), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n812_), .A2(new_n818_), .A3(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1343gat));
  NOR2_X1   g619(.A1(new_n714_), .A2(new_n398_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n780_), .A2(new_n416_), .A3(new_n821_), .A4(new_n782_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n823_));
  OR3_X1    g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n604_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n822_), .B2(new_n604_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n544_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(new_n208_), .ZN(G1344gat));
  AOI22_X1  g626(.A1(new_n824_), .A2(new_n825_), .B1(new_n498_), .B2(new_n496_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(new_n209_), .ZN(G1345gat));
  AOI21_X1  g628(.A(new_n592_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT61), .B(G155gat), .Z(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1346gat));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n825_), .ZN(new_n833_));
  AOI21_X1  g632(.A(G162gat), .B1(new_n833_), .B2(new_n599_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n633_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(G162gat), .B2(new_n835_), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n605_), .A2(new_n416_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n714_), .A3(new_n543_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT123), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n791_), .A2(new_n398_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G169gat), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(KEYINPUT124), .A3(new_n842_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n365_), .A2(new_n605_), .A3(new_n416_), .A4(new_n412_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n791_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n543_), .A3(new_n268_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n842_), .A2(KEYINPUT124), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(KEYINPUT124), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n840_), .A2(G169gat), .A3(new_n848_), .A4(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n847_), .A3(new_n850_), .ZN(G1348gat));
  NAND3_X1  g650(.A1(new_n846_), .A2(new_n269_), .A3(new_n499_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n780_), .A2(new_n782_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n853_), .A2(new_n499_), .A3(new_n844_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n854_), .B2(new_n269_), .ZN(G1349gat));
  NOR3_X1   g654(.A1(new_n845_), .A2(new_n289_), .A3(new_n592_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n701_), .A3(new_n844_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n242_), .ZN(G1350gat));
  OAI21_X1  g657(.A(G190gat), .B1(new_n845_), .B2(new_n633_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n599_), .A2(new_n255_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n845_), .B2(new_n860_), .ZN(G1351gat));
  NAND4_X1  g660(.A1(new_n780_), .A2(new_n821_), .A3(new_n782_), .A4(new_n837_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n543_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n499_), .ZN(new_n866_));
  AND2_X1   g665(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n866_), .B2(new_n867_), .ZN(G1353gat));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n584_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n862_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n701_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT126), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n876_), .A3(new_n701_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n871_), .A2(new_n584_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n875_), .A2(new_n877_), .A3(new_n871_), .A4(new_n584_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1354gat));
  INV_X1    g681(.A(G218gat), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n862_), .A2(new_n883_), .A3(new_n633_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n863_), .A2(new_n599_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(G1355gat));
endmodule


