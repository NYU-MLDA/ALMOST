//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT77), .B(G113gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(G127gat), .A2(G134gat), .ZN(new_n207_));
  INV_X1    g006(.A(G120gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G127gat), .A2(G134gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n206_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n206_), .B1(new_n205_), .B2(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n203_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n206_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n210_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n208_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT78), .A3(new_n211_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT79), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT31), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT31), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(KEYINPUT76), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT72), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT72), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236_));
  INV_X1    g035(.A(G190gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT23), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n227_), .A2(new_n229_), .A3(KEYINPUT24), .A4(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n232_), .A2(new_n241_), .A3(new_n246_), .A4(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n247_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT73), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n226_), .B(new_n255_), .C1(new_n256_), .C2(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT74), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(KEYINPUT22), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n253_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT73), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT74), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n226_), .A4(new_n255_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n251_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n237_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n243_), .A2(KEYINPUT75), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT75), .B1(new_n243_), .B2(new_n245_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n250_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT30), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G43gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(G15gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n272_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G71gat), .B(G99gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(new_n277_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n224_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n280_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n224_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n278_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(G155gat), .B2(G162gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT80), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n292_));
  AND2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n291_), .B(new_n292_), .C1(new_n293_), .C2(new_n287_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n287_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT83), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n293_), .A2(new_n289_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n297_), .A2(KEYINPUT82), .A3(KEYINPUT2), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT81), .B(KEYINPUT2), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n303_), .B(new_n306_), .C1(new_n307_), .C2(new_n297_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n298_), .B(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n302_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n300_), .A2(new_n301_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n301_), .B1(new_n300_), .B2(new_n311_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT29), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G228gat), .ZN(new_n315_));
  INV_X1    g114(.A(G233gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G197gat), .B(G204gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT21), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n319_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n326_), .A2(new_n322_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n321_), .A2(KEYINPUT21), .A3(new_n322_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n314_), .A2(new_n318_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n300_), .A2(new_n311_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT86), .B(KEYINPUT29), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n317_), .B1(new_n334_), .B2(new_n329_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n331_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n286_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n331_), .A2(new_n335_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT28), .ZN(new_n341_));
  INV_X1    g140(.A(new_n286_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n331_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT29), .ZN(new_n345_));
  XOR2_X1   g144(.A(G22gat), .B(G50gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT84), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n345_), .B(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n339_), .A2(new_n344_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n339_), .B2(new_n344_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT90), .B1(new_n270_), .B2(new_n329_), .ZN(new_n355_));
  AOI21_X1  g154(.A(G176gat), .B1(new_n260_), .B2(KEYINPUT73), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n262_), .B1(new_n356_), .B2(new_n255_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n254_), .B1(new_n253_), .B2(new_n259_), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT73), .B1(new_n252_), .B2(G169gat), .ZN(new_n359_));
  NOR4_X1   g158(.A1(new_n358_), .A2(KEYINPUT74), .A3(G176gat), .A4(new_n359_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n247_), .B(new_n269_), .C1(new_n357_), .C2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n249_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n330_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n355_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n246_), .A2(new_n266_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n251_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n256_), .A2(new_n226_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n246_), .A2(KEYINPUT89), .A3(new_n266_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n233_), .A2(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n247_), .A2(new_n373_), .A3(KEYINPUT24), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n247_), .B2(KEYINPUT24), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n230_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n232_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n247_), .A2(KEYINPUT24), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT87), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n247_), .A2(new_n373_), .A3(KEYINPUT24), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n379_), .B(new_n241_), .C1(new_n384_), .C2(new_n230_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n267_), .A2(new_n268_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n329_), .B(new_n371_), .C1(new_n380_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT20), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n354_), .B1(new_n365_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n371_), .B1(new_n380_), .B2(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n330_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n270_), .A2(new_n329_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .A4(new_n354_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT18), .B(G64gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n354_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .A4(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n389_), .B1(new_n355_), .B2(new_n364_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT95), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n411_), .A3(new_n403_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n404_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT96), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n220_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n218_), .A2(new_n211_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n300_), .A3(new_n311_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n220_), .B(KEYINPUT92), .C1(new_n312_), .C2(new_n313_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n417_), .A2(new_n421_), .A3(KEYINPUT4), .A4(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n415_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n423_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n417_), .A2(new_n421_), .A3(new_n424_), .A4(new_n422_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT0), .B(G57gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n414_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n423_), .A2(new_n427_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n429_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n433_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n437_), .A2(KEYINPUT96), .A3(new_n429_), .A4(new_n434_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n413_), .A2(KEYINPUT97), .A3(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT97), .B1(new_n413_), .B2(new_n441_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n401_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n401_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n446_), .B(new_n395_), .C1(new_n407_), .C2(new_n354_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(KEYINPUT91), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n395_), .B1(new_n407_), .B2(new_n354_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n401_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n453_));
  OR3_X1    g252(.A1(new_n428_), .A2(new_n435_), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n417_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n423_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n424_), .B1(new_n415_), .B2(KEYINPUT4), .ZN(new_n457_));
  OAI221_X1 g256(.A(new_n433_), .B1(new_n424_), .B2(new_n455_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n452_), .A2(new_n454_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n352_), .B1(new_n444_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n448_), .A2(new_n451_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n408_), .A2(new_n446_), .ZN(new_n464_));
  AND4_X1   g263(.A1(KEYINPUT98), .A2(new_n464_), .A3(KEYINPUT27), .A4(new_n445_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n449_), .B2(new_n401_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT98), .B1(new_n467_), .B2(new_n464_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n463_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n469_), .A2(new_n441_), .A3(new_n351_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n202_), .B(new_n285_), .C1(new_n461_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n436_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n412_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n411_), .B1(new_n408_), .B2(new_n403_), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n474_), .A2(new_n475_), .B1(new_n397_), .B2(new_n403_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n472_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n413_), .A2(new_n441_), .A3(KEYINPUT97), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n460_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n470_), .B1(new_n479_), .B2(new_n351_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n281_), .A2(new_n284_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT100), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n352_), .A2(new_n469_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n473_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n471_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT6), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT64), .ZN(new_n490_));
  XOR2_X1   g289(.A(G85gat), .B(G92gat), .Z(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  AOI22_X1  g292(.A1(KEYINPUT9), .A2(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n490_), .B(new_n494_), .C1(KEYINPUT9), .C2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT8), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT7), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n490_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n489_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n497_), .B1(new_n502_), .B2(new_n491_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n496_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT66), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n496_), .B(new_n506_), .C1(new_n501_), .C2(new_n503_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n487_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G57gat), .B(G64gat), .Z(new_n509_));
  INV_X1    g308(.A(KEYINPUT11), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G71gat), .A2(G78gat), .ZN(new_n512_));
  INV_X1    g311(.A(G71gat), .ZN(new_n513_));
  INV_X1    g312(.A(G78gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT65), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n509_), .A2(new_n510_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n519_), .A2(new_n504_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n518_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n517_), .B1(new_n510_), .B2(new_n509_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n504_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n487_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .A4(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n519_), .A2(new_n504_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n526_), .ZN(new_n530_));
  OAI211_X1 g329(.A(G230gat), .B(G233gat), .C1(new_n529_), .C2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G204gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT5), .B(G176gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n528_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n528_), .A2(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n535_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n486_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n539_), .A2(new_n486_), .A3(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547_));
  INV_X1    g346(.A(G1gat), .ZN(new_n548_));
  INV_X1    g347(.A(G8gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G1gat), .B(G8gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G29gat), .B(G36gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n553_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT69), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(G229gat), .A3(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n556_), .B(KEYINPUT15), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n553_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n553_), .A2(new_n556_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G197gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT71), .B(G169gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n565_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n546_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n485_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n505_), .A2(new_n507_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n560_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  OAI221_X1 g379(.A(new_n578_), .B1(KEYINPUT35), .B2(new_n580_), .C1(new_n504_), .C2(new_n556_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G190gat), .B(G218gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n588_), .B(new_n589_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n583_), .A2(new_n592_), .A3(new_n584_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT16), .B(G183gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT68), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n553_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n519_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n597_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n576_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n548_), .A3(new_n441_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT38), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n610_), .A2(new_n594_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n576_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n473_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(G1324gat));
  INV_X1    g418(.A(new_n469_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G8gat), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT39), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n613_), .A2(new_n549_), .A3(new_n469_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n617_), .B2(new_n285_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT41), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n613_), .A2(new_n274_), .A3(new_n481_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1326gat));
  OAI21_X1  g428(.A(G22gat), .B1(new_n617_), .B2(new_n351_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n351_), .A2(G22gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n612_), .B2(new_n632_), .ZN(G1327gat));
  INV_X1    g432(.A(new_n594_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n609_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n575_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G29gat), .B1(new_n637_), .B2(new_n441_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n471_), .A2(new_n482_), .A3(KEYINPUT101), .A4(new_n484_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n596_), .B(KEYINPUT102), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n485_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n639_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n485_), .A2(new_n639_), .A3(new_n597_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n574_), .B(new_n610_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n485_), .A2(new_n643_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n640_), .A2(new_n641_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n646_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n654_), .A2(KEYINPUT44), .A3(new_n574_), .A4(new_n610_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n441_), .A2(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n638_), .B1(new_n656_), .B2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n650_), .A2(new_n469_), .A3(new_n655_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(G36gat), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n485_), .A2(new_n662_), .A3(new_n574_), .A4(new_n635_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT103), .B1(new_n663_), .B2(new_n620_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n663_), .A2(KEYINPUT103), .A3(new_n620_), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n661_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n659_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n660_), .B2(G36gat), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n676_), .A2(new_n678_), .A3(KEYINPUT46), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n676_), .B2(KEYINPUT46), .ZN(new_n680_));
  OAI22_X1  g479(.A1(new_n675_), .A2(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1329gat));
  INV_X1    g480(.A(G43gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n637_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(new_n285_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n650_), .A2(G43gat), .A3(new_n481_), .A4(new_n655_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT107), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT107), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT47), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(new_n684_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1330gat));
  NAND2_X1  g491(.A1(new_n656_), .A2(new_n352_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n656_), .A2(KEYINPUT108), .A3(new_n352_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(G50gat), .A3(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n351_), .A2(G50gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n683_), .B2(new_n698_), .ZN(G1331gat));
  NOR2_X1   g498(.A1(new_n545_), .A2(new_n572_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n485_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n611_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n441_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n616_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(G57gat), .A3(new_n441_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n704_), .A2(new_n708_), .ZN(G1332gat));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n469_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G64gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n620_), .A2(G64gat), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT111), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n702_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1333gat));
  NAND3_X1  g515(.A1(new_n702_), .A2(new_n513_), .A3(new_n481_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n707_), .A2(new_n481_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G71gat), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT49), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT49), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT112), .B(new_n717_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1334gat));
  AOI21_X1  g525(.A(new_n514_), .B1(new_n707_), .B2(new_n352_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n702_), .A2(new_n514_), .A3(new_n352_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1335gat));
  NAND2_X1  g529(.A1(new_n701_), .A2(new_n635_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n441_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n609_), .B1(new_n653_), .B2(new_n646_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n700_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n441_), .A2(G85gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1336gat));
  AOI21_X1  g537(.A(G92gat), .B1(new_n732_), .B2(new_n469_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n469_), .A2(G92gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n736_), .B2(new_n740_), .ZN(G1337gat));
  OAI21_X1  g540(.A(G99gat), .B1(new_n735_), .B2(new_n285_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n732_), .A2(new_n492_), .A3(new_n481_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n732_), .A2(new_n493_), .A3(new_n352_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n734_), .A2(new_n352_), .A3(new_n700_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g551(.A(new_n544_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n573_), .B(new_n609_), .C1(new_n753_), .C2(new_n542_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT113), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n545_), .A2(new_n756_), .A3(new_n573_), .A4(new_n609_), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT54), .B(new_n597_), .C1(new_n755_), .C2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n757_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n596_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n758_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n528_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n528_), .B2(new_n763_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n529_), .B1(new_n519_), .B2(new_n508_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n521_), .B1(new_n767_), .B2(new_n527_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n765_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT116), .B1(new_n769_), .B2(new_n536_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  INV_X1    g570(.A(new_n766_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n768_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n528_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n535_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n770_), .A2(new_n771_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT117), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n535_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n770_), .A2(new_n777_), .A3(new_n781_), .A4(new_n771_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n780_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n539_), .A2(new_n572_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT114), .Z(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n539_), .A2(new_n541_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n569_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT118), .Z(new_n789_));
  NAND4_X1  g588(.A1(new_n561_), .A2(G229gat), .A3(G233gat), .A4(new_n563_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n565_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n789_), .A2(new_n790_), .B1(new_n569_), .B2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n787_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n786_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n634_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n771_), .B1(new_n769_), .B2(new_n536_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n780_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n539_), .A3(new_n792_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n803_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n597_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n793_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n797_), .B1(new_n807_), .B2(new_n594_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n799_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n762_), .B1(new_n809_), .B2(new_n610_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n481_), .A2(new_n441_), .A3(new_n483_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT120), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814_), .B2(new_n572_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n610_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n762_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n812_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(KEYINPUT121), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  AOI221_X4 g622(.A(new_n813_), .B1(new_n823_), .B2(new_n821_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n573_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n815_), .B1(new_n826_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g626(.A(new_n208_), .B1(new_n545_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n814_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n208_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n545_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n208_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT122), .B(new_n829_), .C1(new_n830_), .C2(new_n208_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1341gat));
  AOI21_X1  g634(.A(G127gat), .B1(new_n814_), .B2(new_n609_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n822_), .A2(new_n825_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n609_), .A2(G127gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT123), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n836_), .B1(new_n837_), .B2(new_n839_), .ZN(G1342gat));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n821_), .B1(new_n810_), .B2(new_n823_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n814_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n597_), .B1(new_n843_), .B2(new_n824_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G134gat), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n819_), .A2(G134gat), .A3(new_n634_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n841_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT124), .B(new_n846_), .C1(new_n844_), .C2(G134gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1343gat));
  NOR2_X1   g649(.A1(new_n481_), .A2(new_n473_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n818_), .A2(new_n352_), .A3(new_n620_), .A4(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n572_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g656(.A(new_n546_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n854_), .A2(new_n855_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n609_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n609_), .B(new_n860_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1346gat));
  AOI21_X1  g664(.A(G162gat), .B1(new_n861_), .B2(new_n594_), .ZN(new_n866_));
  OAI211_X1 g665(.A(G162gat), .B(new_n641_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1347gat));
  NOR3_X1   g668(.A1(new_n810_), .A2(new_n441_), .A3(new_n285_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n620_), .A2(new_n352_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT126), .B1(new_n872_), .B2(new_n573_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n870_), .A2(new_n874_), .A3(new_n572_), .A4(new_n871_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(G169gat), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n872_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n572_), .A3(new_n256_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n873_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n875_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  NOR2_X1   g681(.A1(new_n872_), .A2(new_n545_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n226_), .ZN(G1349gat));
  NOR2_X1   g683(.A1(new_n872_), .A2(new_n610_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n235_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n265_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n872_), .B2(new_n596_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n594_), .A2(new_n240_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n872_), .B2(new_n889_), .ZN(G1351gat));
  NAND3_X1  g689(.A1(new_n818_), .A2(new_n473_), .A3(new_n469_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n891_), .A2(new_n351_), .A3(new_n481_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n572_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n546_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n609_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  AND2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n897_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n900_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  AOI21_X1  g700(.A(G218gat), .B1(new_n892_), .B2(new_n594_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n597_), .A2(G218gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT127), .Z(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n892_), .B2(new_n904_), .ZN(G1355gat));
endmodule


