//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT7), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n205_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n204_), .A2(new_n205_), .A3(new_n213_), .A4(new_n210_), .ZN(new_n214_));
  OR2_X1    g013(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(KEYINPUT9), .A3(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(KEYINPUT9), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n209_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n212_), .A2(new_n214_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT35), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G232gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT34), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n228_), .A2(new_n231_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n212_), .A2(new_n214_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n220_), .B2(new_n227_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n220_), .A2(new_n227_), .A3(new_n238_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT73), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n231_), .B(KEYINPUT15), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n236_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n235_), .A2(new_n232_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(new_n236_), .B2(KEYINPUT74), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  OAI221_X1 g050(.A(new_n236_), .B1(KEYINPUT74), .B2(new_n249_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G190gat), .B(G218gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G134gat), .B(G162gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT36), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n256_), .A2(KEYINPUT36), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(KEYINPUT75), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT75), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n251_), .A2(new_n252_), .A3(new_n262_), .A4(new_n259_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(KEYINPUT37), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n264_), .A2(KEYINPUT77), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT77), .B1(new_n264_), .B2(new_n266_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G127gat), .B(G155gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT16), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G183gat), .B(G211gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT17), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT78), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G15gat), .B(G22gat), .ZN(new_n277_));
  INV_X1    g076(.A(G1gat), .ZN(new_n278_));
  INV_X1    g077(.A(G8gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT14), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G8gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  NAND2_X1  g082(.A1(G231gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G57gat), .B(G64gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n287_));
  XOR2_X1   g086(.A(G71gat), .B(G78gat), .Z(new_n288_));
  OR2_X1    g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(KEYINPUT11), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n285_), .B(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n273_), .A2(new_n274_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT70), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n276_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n293_), .B1(new_n298_), .B2(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n269_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G230gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT64), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n220_), .A2(new_n227_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n237_), .A2(new_n305_), .A3(new_n292_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT68), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n228_), .A2(new_n308_), .A3(new_n292_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n228_), .A2(new_n292_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n304_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n304_), .B1(new_n228_), .B2(new_n292_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n292_), .A2(KEYINPUT70), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n289_), .B(new_n298_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n314_), .B1(new_n242_), .B2(new_n318_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n228_), .A2(KEYINPUT12), .A3(new_n292_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n313_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n312_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G120gat), .B(G148gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT5), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G176gat), .B(G204gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  OR2_X1    g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n327_), .A2(new_n328_), .B1(new_n331_), .B2(new_n329_), .ZN(new_n332_));
  OR3_X1    g131(.A1(new_n330_), .A2(new_n332_), .A3(KEYINPUT72), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT72), .B1(new_n330_), .B2(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n301_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT79), .ZN(new_n338_));
  XOR2_X1   g137(.A(G8gat), .B(G36gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT18), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT91), .B1(new_n348_), .B2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT91), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(G204gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(G197gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n347_), .B1(new_n354_), .B2(KEYINPUT93), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n354_), .A2(KEYINPUT93), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n349_), .A2(new_n352_), .A3(new_n346_), .A4(new_n353_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n359_), .A2(new_n345_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G197gat), .B(G204gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(new_n346_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(G204gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n353_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n360_), .A2(new_n367_), .A3(KEYINPUT92), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT92), .B1(new_n360_), .B2(new_n367_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n358_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n371_));
  INV_X1    g170(.A(G190gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(KEYINPUT26), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT26), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(KEYINPUT25), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n380_), .A2(G183gat), .B1(new_n372_), .B2(KEYINPUT26), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n376_), .A2(new_n379_), .A3(KEYINPUT84), .A4(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT24), .ZN(new_n387_));
  INV_X1    g186(.A(G169gat), .ZN(new_n388_));
  INV_X1    g187(.A(G176gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n390_), .A2(new_n393_), .A3(KEYINPUT85), .A4(new_n394_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n386_), .A2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n393_), .A2(new_n394_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n377_), .A2(new_n378_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n404_), .B1(G190gat), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G169gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT20), .B1(new_n370_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT92), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT90), .B1(new_n365_), .B2(KEYINPUT21), .ZN(new_n413_));
  AOI211_X1 g212(.A(new_n361_), .B(new_n346_), .C1(new_n364_), .C2(new_n353_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n359_), .A2(new_n345_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n360_), .A2(new_n367_), .A3(KEYINPUT92), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n357_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT25), .B(G183gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT26), .B(G190gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(new_n401_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n395_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n404_), .B1(G183gat), .B2(G190gat), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n423_), .A2(new_n424_), .B1(new_n425_), .B2(new_n408_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n419_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G226gat), .A2(G233gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT19), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n411_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n370_), .B2(new_n410_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n358_), .B(new_n426_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n344_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n429_), .B1(new_n411_), .B2(new_n427_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n343_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G155gat), .B(G162gat), .Z(new_n442_));
  OR3_X1    g241(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(KEYINPUT2), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(KEYINPUT2), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n443_), .B(new_n444_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT1), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n442_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .A4(new_n445_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G127gat), .B(G134gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G120gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n453_), .A2(new_n458_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n464_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n441_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G85gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n453_), .A2(new_n458_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n461_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n453_), .A2(new_n458_), .A3(new_n461_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n441_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n468_), .A2(new_n473_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n473_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(KEYINPUT4), .A3(new_n477_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n440_), .B1(new_n482_), .B2(new_n466_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n483_), .B2(new_n478_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n436_), .A2(new_n439_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n342_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n386_), .A2(new_n402_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n434_), .B(KEYINPUT20), .C1(new_n419_), .C2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(new_n429_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n432_), .B1(new_n419_), .B2(new_n488_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n425_), .A2(new_n408_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n423_), .A2(new_n424_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n370_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n431_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n487_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n437_), .A2(new_n342_), .A3(new_n438_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n437_), .A2(KEYINPUT95), .A3(new_n438_), .A4(new_n342_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n484_), .A2(KEYINPUT33), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n503_), .B(new_n481_), .C1(new_n483_), .C2(new_n478_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n476_), .A2(new_n477_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n440_), .B1(new_n505_), .B2(KEYINPUT97), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n506_), .B1(KEYINPUT97), .B2(new_n505_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n482_), .A2(new_n440_), .A3(new_n466_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n508_), .A2(new_n473_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n502_), .A2(new_n504_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n486_), .B1(new_n501_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n474_), .A2(KEYINPUT29), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n370_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G228gat), .A2(G233gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n370_), .A2(new_n514_), .A3(new_n512_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G78gat), .B(G106gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n474_), .A2(KEYINPUT29), .ZN(new_n523_));
  XOR2_X1   g322(.A(G22gat), .B(G50gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT28), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n523_), .B(new_n525_), .ZN(new_n526_));
  AND4_X1   g325(.A1(KEYINPUT94), .A2(new_n520_), .A3(new_n522_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n529_), .A2(new_n526_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT98), .B1(new_n511_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT98), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n509_), .A2(new_n507_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n468_), .A2(new_n479_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n503_), .B1(new_n536_), .B2(new_n481_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n504_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n500_), .B2(new_n499_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n531_), .B(new_n534_), .C1(new_n540_), .C2(new_n486_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n485_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT27), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n499_), .A2(new_n543_), .A3(new_n500_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n487_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT27), .A3(new_n498_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n532_), .A2(new_n542_), .A3(new_n544_), .A4(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n533_), .A2(new_n541_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(new_n550_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G71gat), .B(G99gat), .ZN(new_n553_));
  INV_X1    g352(.A(G43gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT86), .B(G15gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  MUX2_X1   g358(.A(new_n551_), .B(new_n552_), .S(new_n559_), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n461_), .B(KEYINPUT31), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n561_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n548_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n548_), .A2(KEYINPUT99), .A3(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n544_), .A2(new_n546_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(new_n532_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n565_), .A2(new_n485_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n568_), .A2(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT81), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n283_), .A2(new_n231_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT80), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n283_), .A2(new_n231_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n283_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n244_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n580_), .A3(new_n575_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n582_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n582_), .B2(new_n585_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n574_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n582_), .A2(new_n585_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n588_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(KEYINPUT81), .A3(new_n589_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n573_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n338_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n485_), .B(KEYINPUT100), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n278_), .A3(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n258_), .A2(new_n260_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n573_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n300_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n336_), .A2(new_n605_), .A3(new_n597_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(new_n485_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n602_), .B1(new_n278_), .B2(new_n608_), .ZN(new_n609_));
  MUX2_X1   g408(.A(new_n602_), .B(new_n609_), .S(KEYINPUT38), .Z(G1324gat));
  AOI21_X1  g409(.A(new_n279_), .B1(new_n607_), .B2(new_n570_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT39), .Z(new_n612_));
  NAND3_X1  g411(.A1(new_n599_), .A2(new_n279_), .A3(new_n570_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(KEYINPUT40), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1325gat));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n607_), .B2(new_n564_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT41), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n599_), .A2(new_n619_), .A3(new_n564_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1326gat));
  INV_X1    g422(.A(G22gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n607_), .B2(new_n532_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT42), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n599_), .A2(new_n624_), .A3(new_n532_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1327gat));
  OAI21_X1  g427(.A(KEYINPUT43), .B1(new_n573_), .B2(new_n269_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n572_), .A2(new_n571_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n548_), .A2(KEYINPUT99), .A3(new_n565_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT99), .B1(new_n548_), .B2(new_n565_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n267_), .A2(new_n268_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n629_), .A2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n336_), .A2(new_n300_), .A3(new_n597_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n600_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n603_), .A2(new_n605_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT101), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n336_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n598_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n542_), .A2(G29gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT102), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n644_), .B1(new_n648_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(new_n570_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G36gat), .B1(new_n643_), .B2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n652_), .A2(G36gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT103), .B1(new_n648_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT45), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n648_), .A2(KEYINPUT103), .A3(new_n654_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n662_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n653_), .A2(new_n664_), .A3(new_n659_), .A4(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1329gat));
  OAI21_X1  g465(.A(new_n554_), .B1(new_n648_), .B2(new_n565_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n564_), .A2(G43gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n643_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n669_), .B(new_n670_), .Z(G1330gat));
  OR3_X1    g470(.A1(new_n648_), .A2(G50gat), .A3(new_n531_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n641_), .A2(new_n532_), .A3(new_n642_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT106), .A3(G50gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT106), .B1(new_n673_), .B2(G50gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n301_), .A2(new_n335_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT107), .Z(new_n678_));
  INV_X1    g477(.A(new_n597_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n573_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(G57gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(new_n601_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n335_), .A2(new_n605_), .A3(new_n679_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n604_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n542_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n682_), .A2(new_n686_), .ZN(G1332gat));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n684_), .B2(new_n570_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT48), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n680_), .A2(new_n688_), .A3(new_n570_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1333gat));
  INV_X1    g491(.A(G71gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n680_), .A2(new_n693_), .A3(new_n564_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n684_), .B2(new_n564_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT109), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(G1334gat));
  NOR2_X1   g499(.A1(new_n531_), .A2(G78gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n680_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G78gat), .B1(new_n685_), .B2(new_n531_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT50), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT50), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(G1335gat));
  NOR3_X1   g506(.A1(new_n335_), .A2(new_n300_), .A3(new_n679_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n629_), .B2(new_n636_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711_), .B2(new_n542_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n646_), .A2(new_n335_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n633_), .A2(new_n597_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT111), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n633_), .A2(new_n716_), .A3(new_n597_), .A4(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n221_), .A3(new_n601_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n712_), .A2(new_n719_), .ZN(G1336gat));
  OAI21_X1  g519(.A(G92gat), .B1(new_n711_), .B2(new_n652_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n222_), .A3(new_n570_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1337gat));
  AND3_X1   g522(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n634_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n564_), .B(new_n708_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G99gat), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n215_), .A2(new_n217_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n565_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n718_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n728_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n726_), .A2(G99gat), .B1(new_n718_), .B2(new_n730_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .A3(new_n728_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n735_), .B2(new_n728_), .ZN(new_n739_));
  INV_X1    g538(.A(G99gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n710_), .B2(new_n564_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n729_), .B(new_n565_), .C1(new_n715_), .C2(new_n717_), .ZN(new_n742_));
  OAI211_X1 g541(.A(KEYINPUT112), .B(KEYINPUT51), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n739_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n737_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n737_), .A2(new_n744_), .A3(KEYINPUT114), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1338gat));
  NAND3_X1  g548(.A1(new_n718_), .A2(new_n216_), .A3(new_n532_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n710_), .A2(new_n532_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G106gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT52), .B(new_n216_), .C1(new_n710_), .C2(new_n532_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT53), .ZN(G1339gat));
  AND3_X1   g555(.A1(new_n592_), .A2(new_n596_), .A3(new_n300_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT115), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n757_), .C1(new_n330_), .C2(new_n332_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n762_), .B(new_n763_), .C1(new_n268_), .C2(new_n267_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n269_), .B2(new_n762_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n327_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n597_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n237_), .A2(new_n305_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n292_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n314_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n241_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n239_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n317_), .B1(new_n776_), .B2(new_n237_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n777_), .B2(new_n314_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n771_), .B1(new_n778_), .B2(new_n313_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT118), .B1(new_n778_), .B2(new_n313_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n770_), .A2(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n321_), .A2(KEYINPUT116), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT118), .A3(KEYINPUT55), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n319_), .A2(new_n320_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT117), .B1(new_n785_), .B2(new_n310_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n778_), .A2(new_n787_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n304_), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(new_n784_), .A3(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n326_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n326_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n769_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n327_), .A2(new_n328_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n580_), .B1(new_n283_), .B2(new_n231_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n588_), .B1(new_n584_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n579_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n581_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n589_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n603_), .B1(new_n793_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT57), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n327_), .A2(new_n589_), .A3(new_n798_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT58), .B(new_n802_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT120), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n790_), .A2(new_n326_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n326_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(KEYINPUT58), .A4(new_n802_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n802_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n635_), .A2(new_n804_), .A3(new_n811_), .A4(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n800_), .B2(KEYINPUT119), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n818_), .B(new_n603_), .C1(new_n793_), .C2(new_n799_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n801_), .B(new_n815_), .C1(new_n817_), .C2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n767_), .B1(new_n605_), .B2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n565_), .A2(new_n600_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n571_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n679_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n815_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n828_), .A2(KEYINPUT121), .B1(KEYINPUT57), .B2(new_n800_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n815_), .C1(new_n817_), .C2(new_n819_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n300_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n827_), .B1(new_n832_), .B2(new_n767_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n823_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n679_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n826_), .B1(new_n837_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n335_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n824_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n835_), .A2(new_n336_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n839_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n824_), .B2(new_n300_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n300_), .A2(G127gat), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT122), .Z(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n835_), .B2(new_n847_), .ZN(G1342gat));
  NAND2_X1  g647(.A1(new_n828_), .A2(KEYINPUT121), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n801_), .A3(new_n831_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n767_), .B1(new_n850_), .B2(new_n605_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n827_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n635_), .B(new_n834_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G134gat), .ZN(new_n854_));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n824_), .A2(new_n855_), .A3(new_n603_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n854_), .A2(KEYINPUT123), .A3(new_n856_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1343gat));
  OR2_X1    g660(.A1(new_n765_), .A2(new_n766_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n820_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n300_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n564_), .A2(new_n531_), .ZN(new_n865_));
  AND4_X1   g664(.A1(new_n652_), .A2(new_n864_), .A3(new_n601_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n679_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n336_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n873_), .A3(new_n300_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n866_), .B2(new_n300_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n872_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n876_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n874_), .A3(new_n871_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n866_), .B2(new_n603_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n635_), .A2(G162gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n866_), .B2(new_n883_), .ZN(G1347gat));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n851_), .A2(new_n532_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n565_), .A2(new_n652_), .A3(new_n601_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n679_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n885_), .B1(new_n888_), .B2(G169gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n531_), .B(new_n887_), .C1(new_n832_), .C2(new_n767_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n885_), .B(G169gat), .C1(new_n890_), .C2(new_n597_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT22), .B(G169gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n679_), .A2(new_n893_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT126), .Z(new_n895_));
  OAI22_X1  g694(.A1(new_n889_), .A2(new_n892_), .B1(new_n890_), .B2(new_n895_), .ZN(G1348gat));
  NAND3_X1  g695(.A1(new_n886_), .A2(new_n336_), .A3(new_n887_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n821_), .A2(new_n532_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n336_), .A2(G176gat), .A3(new_n887_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n389_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NAND2_X1  g699(.A1(new_n887_), .A2(new_n300_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n405_), .B1(new_n898_), .B2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n420_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n886_), .B2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n890_), .B2(new_n269_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n603_), .A2(new_n421_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n890_), .B2(new_n907_), .ZN(G1351gat));
  NOR2_X1   g707(.A1(new_n652_), .A2(new_n485_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n864_), .A2(new_n865_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n679_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n336_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g713(.A(new_n605_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n910_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n916_), .B(new_n917_), .Z(G1354gat));
  AND2_X1   g717(.A1(new_n910_), .A2(new_n603_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G218gat), .B1(new_n919_), .B2(new_n920_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n635_), .A2(G218gat), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n922_), .B1(new_n910_), .B2(new_n923_), .ZN(G1355gat));
endmodule


