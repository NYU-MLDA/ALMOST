//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT8), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT65), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n207_), .B(new_n209_), .C1(new_n215_), .C2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n218_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n204_), .A2(KEYINPUT9), .A3(new_n205_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n214_), .A2(new_n225_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n221_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n206_), .B1(new_n229_), .B2(new_n214_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n222_), .B(new_n228_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G43gat), .B(G50gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G36gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G29gat), .ZN(new_n237_));
  INV_X1    g036(.A(G29gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G36gat), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n237_), .A2(new_n239_), .A3(KEYINPUT69), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT69), .B1(new_n237_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n235_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n238_), .A2(G36gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n236_), .A2(G29gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n237_), .A2(new_n239_), .A3(KEYINPUT69), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n234_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT70), .B1(new_n233_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n207_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n225_), .A2(new_n226_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n214_), .A2(new_n227_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n251_), .A2(new_n231_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .A4(new_n222_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT34), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT71), .B1(new_n260_), .B2(KEYINPUT35), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT15), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n249_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n242_), .A2(new_n248_), .A3(KEYINPUT15), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n265_), .B2(new_n233_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(KEYINPUT35), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G134gat), .B(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT36), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n258_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n258_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n268_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT73), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(new_n281_), .A3(new_n275_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n273_), .B(KEYINPUT36), .Z(new_n284_));
  AOI21_X1  g083(.A(new_n277_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n284_), .ZN(new_n286_));
  AOI211_X1 g085(.A(KEYINPUT74), .B(new_n286_), .C1(new_n280_), .C2(new_n282_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n276_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT37), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n276_), .A2(KEYINPUT72), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n284_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(new_n276_), .A3(KEYINPUT72), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G127gat), .B(G155gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(G183gat), .B(G211gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  XNOR2_X1  g110(.A(G57gat), .B(G64gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT11), .ZN(new_n313_));
  XOR2_X1   g112(.A(G71gat), .B(G78gat), .Z(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n314_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n312_), .A2(KEYINPUT11), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n311_), .B(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n302_), .B1(new_n319_), .B2(KEYINPUT17), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(KEYINPUT17), .B2(new_n302_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT76), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n297_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G8gat), .B(G36gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT19), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338_));
  OR2_X1    g137(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n337_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G169gat), .ZN(new_n344_));
  INV_X1    g143(.A(G176gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(KEYINPUT80), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(G169gat), .B2(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT24), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT23), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n346_), .A2(new_n348_), .A3(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n343_), .A2(new_n351_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n339_), .A2(new_n340_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(G190gat), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(G176gat), .B1(KEYINPUT81), .B2(KEYINPUT22), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G169gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G197gat), .B(G204gat), .Z(new_n363_));
  INV_X1    g162(.A(KEYINPUT21), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(KEYINPUT91), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n363_), .A2(KEYINPUT21), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT100), .B1(new_n362_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n362_), .A2(new_n373_), .A3(KEYINPUT100), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n353_), .B1(G183gat), .B2(G190gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n350_), .B(KEYINPUT99), .Z(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT22), .B(G169gat), .Z(new_n380_));
  OAI211_X1 g179(.A(new_n378_), .B(new_n379_), .C1(G176gat), .C2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT97), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n337_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n337_), .A2(new_n382_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT25), .B(G183gat), .Z(new_n385_));
  NOR3_X1   g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT98), .B(KEYINPUT24), .Z(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n388_), .B(new_n353_), .C1(new_n349_), .C2(new_n387_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n381_), .B(new_n372_), .C1(new_n386_), .C2(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(KEYINPUT20), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n336_), .B1(new_n377_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n372_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n381_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n373_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT96), .B1(new_n393_), .B2(KEYINPUT20), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n397_), .A2(new_n335_), .A3(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n333_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT104), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n335_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n376_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n391_), .B(new_n336_), .C1(new_n403_), .C2(new_n374_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n404_), .A3(new_n332_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT27), .A4(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT27), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n402_), .A2(new_n404_), .A3(new_n332_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n332_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n400_), .A2(KEYINPUT27), .A3(new_n405_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT104), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT90), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n373_), .B2(KEYINPUT92), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G141gat), .A2(G148gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G141gat), .A2(G148gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(KEYINPUT1), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(KEYINPUT1), .ZN(new_n424_));
  AOI211_X1 g223(.A(new_n418_), .B(new_n420_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n426_));
  NOR2_X1   g225(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n428_), .B(KEYINPUT86), .C1(new_n430_), .C2(new_n431_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n418_), .B2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(KEYINPUT88), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT2), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n420_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n419_), .B1(new_n442_), .B2(KEYINPUT88), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n441_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n436_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G155gat), .B(G162gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT89), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n425_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT29), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n417_), .B1(new_n456_), .B2(new_n372_), .ZN(new_n457_));
  OAI221_X1 g256(.A(new_n373_), .B1(KEYINPUT92), .B2(new_n416_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT93), .Z(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT28), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n454_), .A2(new_n464_), .A3(new_n455_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n425_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n448_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n452_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT28), .B1(new_n468_), .B2(KEYINPUT29), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G22gat), .B(G50gat), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n465_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT94), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n462_), .B1(new_n463_), .B2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n471_), .A2(new_n472_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(KEYINPUT94), .A3(new_n459_), .A4(new_n461_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n457_), .A2(new_n458_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n460_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n474_), .A2(new_n476_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT31), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G43gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G227gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(G15gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n489_), .B(new_n492_), .Z(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G127gat), .B(G134gat), .Z(new_n495_));
  INV_X1    g294(.A(G120gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G113gat), .ZN(new_n497_));
  INV_X1    g296(.A(G113gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G120gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G127gat), .B(G134gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT83), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n495_), .B2(new_n500_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n494_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n494_), .A2(new_n507_), .ZN(new_n509_));
  OR3_X1    g308(.A1(new_n486_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n468_), .A2(new_n511_), .A3(new_n507_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n452_), .B1(new_n436_), .B2(new_n449_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n507_), .B1(new_n516_), .B2(new_n425_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT102), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n501_), .A2(new_n518_), .A3(new_n503_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n521_), .B(new_n466_), .C1(new_n467_), .C2(new_n452_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n522_), .A3(KEYINPUT4), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n517_), .A2(new_n522_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n515_), .A2(new_n523_), .B1(new_n524_), .B2(new_n513_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G1gat), .B(G29gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n202_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT0), .B(G57gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n517_), .A2(new_n522_), .A3(new_n513_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n517_), .A2(KEYINPUT4), .A3(new_n522_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n512_), .A2(new_n514_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n531_), .B(new_n529_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n486_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n510_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n414_), .A2(new_n482_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT103), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n529_), .A2(KEYINPUT33), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n531_), .B(new_n543_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n529_), .B1(new_n524_), .B2(new_n514_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n523_), .A2(new_n513_), .A3(new_n512_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n402_), .A2(new_n404_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n333_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n405_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n540_), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n408_), .A2(new_n409_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n525_), .A2(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT103), .A4(new_n542_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n557_), .B(new_n558_), .C1(new_n535_), .C2(new_n530_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n555_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n474_), .A2(new_n476_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n479_), .A2(new_n481_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n482_), .A2(new_n411_), .A3(new_n536_), .A4(new_n413_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n510_), .A2(new_n537_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n539_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G169gat), .B(G197gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n309_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n265_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT78), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n309_), .B2(new_n255_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n309_), .B(new_n255_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n577_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n571_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(new_n581_), .A3(new_n571_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n233_), .B(new_n318_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT64), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT66), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n233_), .A2(new_n594_), .A3(new_n318_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n589_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G120gat), .B(G148gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n593_), .A2(new_n597_), .A3(new_n603_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n605_), .A2(KEYINPUT68), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT68), .B1(new_n605_), .B2(new_n606_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT13), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT13), .B1(new_n607_), .B2(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n568_), .A2(new_n586_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n327_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n536_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n304_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  INV_X1    g417(.A(new_n288_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n568_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n324_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n613_), .A2(new_n621_), .A3(new_n586_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n304_), .B1(new_n623_), .B2(new_n616_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT105), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT107), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n620_), .A2(new_n414_), .A3(new_n622_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT106), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(G8gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n629_), .B2(G8gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(KEYINPUT107), .A3(new_n631_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n634_), .A2(new_n636_), .A3(KEYINPUT39), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n628_), .B(new_n638_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n615_), .A2(new_n305_), .A3(new_n414_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n627_), .B1(new_n637_), .B2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(new_n636_), .A3(KEYINPUT39), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT40), .A3(new_n639_), .A4(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1325gat));
  INV_X1    g444(.A(new_n567_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n491_), .B1(new_n623_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT41), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n615_), .A2(new_n491_), .A3(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1326gat));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n615_), .A2(new_n651_), .A3(new_n482_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n623_), .A2(new_n482_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(G22gat), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT42), .B(new_n651_), .C1(new_n623_), .C2(new_n482_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT108), .ZN(G1327gat));
  AOI21_X1  g457(.A(new_n646_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT109), .B(new_n294_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n659_), .A2(new_n539_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT43), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT43), .B1(new_n290_), .B2(new_n295_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n659_), .B2(new_n539_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT110), .B(new_n665_), .C1(new_n659_), .C2(new_n539_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n613_), .A2(new_n324_), .A3(new_n586_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(KEYINPUT43), .A2(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n669_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(new_n238_), .A3(new_n536_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n324_), .A2(new_n288_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n614_), .A2(new_n616_), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n238_), .B2(new_n680_), .ZN(G1328gat));
  OAI211_X1 g480(.A(new_n672_), .B(new_n414_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n414_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n614_), .A2(new_n679_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n683_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT46), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n688_), .B1(new_n682_), .B2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n693_), .A2(KEYINPUT112), .A3(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1329gat));
  NAND2_X1  g495(.A1(new_n646_), .A2(G43gat), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n677_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n614_), .A2(new_n646_), .A3(new_n679_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n488_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n698_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1330gat));
  INV_X1    g503(.A(G50gat), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n677_), .A2(new_n705_), .A3(new_n563_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n614_), .A2(new_n482_), .A3(new_n679_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(new_n707_), .ZN(G1331gat));
  INV_X1    g507(.A(new_n613_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(new_n621_), .A3(new_n585_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n620_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n536_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n568_), .A2(new_n709_), .A3(new_n585_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n327_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n536_), .B1(new_n715_), .B2(KEYINPUT114), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(KEYINPUT114), .B2(new_n715_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n717_), .B2(new_n712_), .ZN(G1332gat));
  OAI21_X1  g517(.A(G64gat), .B1(new_n711_), .B2(new_n684_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT48), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n684_), .A2(G64gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n715_), .B2(new_n721_), .ZN(G1333gat));
  NAND3_X1  g521(.A1(new_n710_), .A2(new_n620_), .A3(new_n646_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(G71gat), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G71gat), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n567_), .A2(G71gat), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n725_), .A2(new_n726_), .B1(new_n715_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT116), .Z(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n711_), .B2(new_n563_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT50), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n563_), .A2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n715_), .B2(new_n732_), .ZN(G1335gat));
  AND2_X1   g532(.A1(new_n714_), .A2(new_n679_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n202_), .A3(new_n616_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n670_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n709_), .A2(new_n324_), .A3(new_n585_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n736_), .A2(new_n536_), .A3(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n739_), .B2(new_n202_), .ZN(G1336gat));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n203_), .A3(new_n414_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n736_), .A2(new_n684_), .A3(new_n738_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n203_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n670_), .A2(new_n646_), .A3(new_n737_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G99gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n734_), .A2(new_n646_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n748_), .B(new_n749_), .Z(G1338gat));
  NAND3_X1  g549(.A1(new_n734_), .A2(new_n218_), .A3(new_n482_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n670_), .A2(new_n482_), .A3(new_n737_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g556(.A1(new_n414_), .A2(new_n482_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n616_), .A3(new_n646_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n575_), .B(new_n577_), .C1(new_n249_), .C2(new_n572_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n571_), .B1(new_n580_), .B2(new_n576_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(new_n584_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT55), .B1(new_n596_), .B2(new_n589_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n597_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n596_), .A2(KEYINPUT55), .A3(new_n589_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n604_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n604_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n584_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n606_), .B1(new_n773_), .B2(new_n582_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n768_), .B2(KEYINPUT118), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n609_), .A2(new_n763_), .B1(new_n772_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT120), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .A4(new_n619_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n775_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n605_), .A2(new_n606_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT68), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n605_), .A2(KEYINPUT68), .A3(new_n606_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(new_n763_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n619_), .B1(new_n780_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT120), .B1(new_n786_), .B2(KEYINPUT57), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n779_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n778_), .B1(new_n776_), .B2(new_n619_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n606_), .A2(new_n762_), .A3(new_n584_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n771_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n768_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT58), .B(new_n790_), .C1(new_n791_), .C2(new_n768_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n296_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n794_), .A2(new_n296_), .A3(KEYINPUT119), .A4(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n789_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n621_), .B1(new_n788_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n611_), .A2(new_n612_), .A3(new_n586_), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n325_), .A2(new_n802_), .A3(KEYINPUT54), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT54), .B1(new_n325_), .B2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n759_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G113gat), .B1(new_n806_), .B2(new_n585_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  INV_X1    g607(.A(new_n759_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n780_), .A2(new_n785_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n288_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n777_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n786_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n789_), .A2(new_n796_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n324_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n803_), .A2(new_n804_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n808_), .B(new_n809_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n806_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(KEYINPUT59), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n498_), .B1(new_n585_), .B2(KEYINPUT121), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(KEYINPUT121), .B2(new_n498_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n807_), .B1(new_n821_), .B2(new_n823_), .ZN(G1340gat));
  OAI21_X1  g623(.A(new_n496_), .B1(new_n709_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n806_), .B(new_n825_), .C1(KEYINPUT60), .C2(new_n496_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n818_), .B(new_n613_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n828_), .B2(new_n496_), .ZN(G1341gat));
  NAND2_X1  g628(.A1(new_n806_), .A2(new_n324_), .ZN(new_n830_));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n621_), .A2(new_n831_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n818_), .B(new_n833_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT122), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT122), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n806_), .A2(new_n840_), .A3(new_n619_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n818_), .B(new_n296_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n840_), .ZN(G1343gat));
  NAND2_X1  g643(.A1(new_n482_), .A2(new_n567_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n414_), .A2(new_n536_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n800_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n324_), .B1(new_n848_), .B2(new_n814_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n846_), .B(new_n847_), .C1(new_n849_), .C2(new_n817_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n585_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n613_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n850_), .B2(new_n621_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n845_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n858_), .A2(KEYINPUT123), .A3(new_n324_), .A4(new_n847_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n857_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1346gat));
  AOI21_X1  g662(.A(G162gat), .B1(new_n851_), .B2(new_n619_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G162gat), .B1(new_n661_), .B2(new_n662_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT124), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n851_), .B2(new_n866_), .ZN(G1347gat));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n684_), .A2(new_n538_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n563_), .A3(new_n585_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n380_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n874_), .B(new_n871_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT62), .B1(new_n872_), .B2(G169gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n868_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n877_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n879_), .A2(KEYINPUT125), .A3(new_n875_), .A4(new_n873_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1348gat));
  NOR2_X1   g680(.A1(new_n816_), .A2(new_n817_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n869_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n882_), .A2(new_n482_), .A3(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G176gat), .B1(new_n884_), .B2(new_n613_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n482_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n709_), .A2(new_n345_), .A3(new_n883_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  AND2_X1   g687(.A1(new_n324_), .A2(new_n385_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n324_), .A3(new_n869_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n357_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n884_), .A2(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n884_), .A2(new_n296_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G190gat), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n288_), .A2(new_n384_), .A3(new_n383_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n884_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1351gat));
  NOR2_X1   g696(.A1(new_n684_), .A2(new_n616_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n858_), .A2(new_n585_), .A3(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g699(.A1(new_n858_), .A2(new_n613_), .A3(new_n898_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g701(.A1(new_n858_), .A2(new_n898_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n324_), .A2(new_n904_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT126), .Z(new_n906_));
  NOR2_X1   g705(.A1(new_n903_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1354gat));
  OAI21_X1  g708(.A(G218gat), .B1(new_n903_), .B2(new_n297_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n288_), .A2(G218gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n903_), .B2(new_n911_), .ZN(G1355gat));
endmodule


