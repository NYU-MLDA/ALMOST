//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  NOR2_X1   g000(.A1(G197gat), .A2(G204gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT86), .B(G197gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(G204gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT87), .ZN(new_n205_));
  XOR2_X1   g004(.A(G211gat), .B(G218gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(KEYINPUT87), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n205_), .A2(KEYINPUT21), .A3(new_n206_), .A4(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n203_), .A2(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(G197gat), .B2(G204gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n206_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT21), .B2(new_n204_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT26), .B(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT82), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT23), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n222_), .A2(KEYINPUT92), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT92), .B1(new_n222_), .B2(new_n224_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(new_n220_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n219_), .A3(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n208_), .A2(new_n213_), .A3(new_n227_), .A4(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n233_), .A2(KEYINPUT20), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G226gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n208_), .A2(new_n213_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n241_), .A2(new_n222_), .A3(new_n216_), .A4(new_n220_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n229_), .A2(KEYINPUT83), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT83), .B1(new_n244_), .B2(KEYINPUT22), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(new_n230_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n228_), .B(new_n219_), .C1(new_n243_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n234_), .A2(new_n235_), .A3(new_n239_), .A4(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n233_), .A3(KEYINPUT20), .A4(new_n239_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT93), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n240_), .A2(new_n248_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n227_), .A2(new_n232_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n240_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n239_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n252_), .B2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G8gat), .B(G36gat), .Z(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n250_), .B(new_n263_), .C1(new_n252_), .C2(new_n257_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n256_), .A2(new_n239_), .A3(new_n253_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n239_), .B1(new_n234_), .B2(new_n249_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n263_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(KEYINPUT27), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT3), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT2), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G155gat), .B(G162gat), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n283_), .B1(KEYINPUT1), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(KEYINPUT1), .B2(new_n284_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n276_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(new_n278_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n240_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G228gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G78gat), .B(G106gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT90), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n290_), .A2(KEYINPUT29), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G22gat), .B(G50gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(KEYINPUT90), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT88), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n294_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n294_), .A2(new_n306_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n295_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT89), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n311_), .B(new_n295_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n294_), .A2(new_n296_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n303_), .B1(new_n315_), .B2(new_n297_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n275_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G71gat), .B(G99gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G43gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n248_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(G15gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT30), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT31), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n328_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(new_n327_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n328_), .A2(new_n338_), .A3(new_n336_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT96), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n280_), .A2(new_n281_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n332_), .A2(new_n334_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(KEYINPUT95), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT95), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n341_), .B(new_n342_), .C1(new_n344_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n335_), .A2(new_n345_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n346_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n290_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT96), .B1(new_n342_), .B2(new_n343_), .ZN(new_n351_));
  OAI211_X1 g150(.A(KEYINPUT4), .B(new_n347_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n290_), .A2(new_n335_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  OAI21_X1  g162(.A(new_n342_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n353_), .A3(KEYINPUT96), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n358_), .B1(new_n365_), .B2(new_n347_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n359_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n363_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n357_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n340_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n318_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n359_), .A2(KEYINPUT33), .A3(new_n363_), .A4(new_n367_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT97), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n347_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n363_), .B1(new_n378_), .B2(new_n358_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n358_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT98), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n356_), .A2(new_n357_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT98), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n379_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n368_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n386_), .A2(new_n388_), .A3(new_n265_), .A4(new_n266_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT99), .B1(new_n377_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT97), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n376_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT99), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n382_), .A2(new_n385_), .B1(new_n368_), .B2(new_n387_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n392_), .A2(new_n267_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n258_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT32), .B(new_n264_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n372_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT100), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n372_), .A2(new_n398_), .A3(KEYINPUT100), .A4(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(KEYINPUT101), .A3(new_n317_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n373_), .B1(new_n313_), .B2(new_n316_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n274_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT101), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n404_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n313_), .A2(new_n316_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n340_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n375_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G29gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G43gat), .B(G50gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G1gat), .B(G8gat), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G1gat), .A2(G8gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT14), .ZN(new_n424_));
  INV_X1    g223(.A(G22gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n323_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G15gat), .A2(G22gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(KEYINPUT77), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(KEYINPUT77), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n422_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(new_n421_), .A3(new_n433_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n420_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n420_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n436_), .A2(new_n438_), .A3(KEYINPUT79), .A4(new_n420_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G229gat), .A2(G233gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n442_), .A2(new_n443_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n436_), .A2(new_n438_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n420_), .B(KEYINPUT15), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n449_), .B(new_n445_), .C1(new_n450_), .C2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT80), .B1(new_n444_), .B2(new_n445_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n448_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G113gat), .B(G141gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT81), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G169gat), .B(G197gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n448_), .A2(new_n453_), .A3(new_n454_), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n417_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G85gat), .ZN(new_n466_));
  INV_X1    g265(.A(G92gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT9), .B1(new_n471_), .B2(KEYINPUT66), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  AND4_X1   g272(.A1(KEYINPUT66), .A2(new_n468_), .A3(KEYINPUT9), .A4(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n468_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT67), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT68), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT68), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n484_));
  INV_X1    g283(.A(G99gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT65), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n486_), .A2(KEYINPUT65), .A3(new_n487_), .A4(new_n488_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n483_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n468_), .A2(KEYINPUT66), .A3(new_n473_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT9), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n471_), .A2(KEYINPUT66), .A3(KEYINPUT9), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n468_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n476_), .A2(new_n494_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n478_), .A2(new_n480_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT68), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT68), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT8), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n471_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n478_), .A2(new_n480_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n506_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT69), .B(new_n471_), .C1(new_n514_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT8), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n509_), .A2(new_n503_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT69), .B1(new_n520_), .B2(new_n471_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n513_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n502_), .A2(new_n522_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT70), .Z(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n502_), .B2(new_n522_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT71), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G230gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT64), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT72), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(KEYINPUT73), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n500_), .B1(new_n499_), .B2(new_n468_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n483_), .A2(new_n493_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n471_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT8), .A3(new_n518_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n544_), .A2(new_n501_), .B1(new_n548_), .B2(new_n513_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n541_), .B1(new_n549_), .B2(new_n529_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n536_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n502_), .A2(new_n522_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n529_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n550_), .A2(new_n551_), .A3(new_n530_), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n534_), .A2(new_n558_), .A3(new_n536_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n538_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G120gat), .B(G148gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT5), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n560_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n529_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n450_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(KEYINPUT17), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n572_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n549_), .A2(new_n420_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT34), .Z(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT74), .Z(new_n587_));
  OAI211_X1 g386(.A(new_n582_), .B(new_n587_), .C1(new_n452_), .C2(new_n549_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT75), .B1(new_n549_), .B2(new_n452_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n584_), .A2(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n588_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT76), .ZN(new_n595_));
  XOR2_X1   g394(.A(G134gat), .B(G162gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n593_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n592_), .A2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n598_), .A2(KEYINPUT37), .A3(new_n600_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n569_), .A2(new_n581_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n465_), .A2(new_n606_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n607_), .A2(G1gat), .A3(new_n373_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT38), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n417_), .A2(new_n601_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n569_), .A2(new_n464_), .A3(new_n581_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n373_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n609_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  NOR3_X1   g415(.A1(new_n607_), .A2(G8gat), .A3(new_n275_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G8gat), .B1(new_n613_), .B2(new_n275_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(KEYINPUT39), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(KEYINPUT39), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(G1325gat));
  OAI21_X1  g422(.A(G15gat), .B1(new_n613_), .B2(new_n416_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT41), .Z(new_n625_));
  INV_X1    g424(.A(new_n607_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n323_), .A3(new_n340_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(G1326gat));
  OAI21_X1  g427(.A(G22gat), .B1(new_n613_), .B2(new_n317_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT42), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n425_), .A3(new_n413_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1327gat));
  NAND2_X1  g431(.A1(new_n601_), .A2(new_n581_), .ZN(new_n633_));
  NOR4_X1   g432(.A1(new_n417_), .A2(new_n464_), .A3(new_n569_), .A4(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n372_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT104), .B1(new_n636_), .B2(KEYINPUT105), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n415_), .A2(new_n416_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n375_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n641_), .B2(new_n605_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n605_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n417_), .A2(KEYINPUT43), .A3(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n569_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n463_), .A3(new_n581_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n637_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n406_), .A2(new_n317_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n409_), .B1(new_n649_), .B2(new_n411_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n340_), .B1(new_n650_), .B2(new_n407_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n638_), .B(new_n605_), .C1(new_n651_), .C2(new_n375_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n417_), .B2(new_n643_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n647_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT105), .B1(new_n654_), .B2(KEYINPUT104), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n648_), .B1(new_n655_), .B2(KEYINPUT44), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n372_), .A2(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n635_), .B1(new_n656_), .B2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659_));
  INV_X1    g458(.A(G36gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n656_), .B2(new_n274_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n634_), .A2(new_n660_), .A3(new_n274_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT45), .Z(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n663_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n666_));
  AOI211_X1 g465(.A(new_n666_), .B(new_n647_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n636_), .B1(new_n667_), .B2(KEYINPUT105), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n275_), .B1(new_n668_), .B2(new_n648_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n665_), .B(KEYINPUT46), .C1(new_n669_), .C2(new_n660_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(new_n670_), .ZN(G1329gat));
  INV_X1    g470(.A(KEYINPUT47), .ZN(new_n672_));
  INV_X1    g471(.A(G43gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n656_), .B2(new_n340_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n634_), .A2(new_n673_), .A3(new_n340_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n416_), .B1(new_n668_), .B2(new_n648_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT47), .B(new_n675_), .C1(new_n678_), .C2(new_n673_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n634_), .B2(new_n413_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n413_), .A2(G50gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n656_), .B2(new_n682_), .ZN(G1331gat));
  NOR2_X1   g482(.A1(new_n605_), .A2(new_n581_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n569_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT106), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n417_), .A2(new_n463_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n372_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n646_), .A2(new_n463_), .A3(new_n581_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n611_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(new_n372_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n693_), .B2(new_n689_), .ZN(G1332gat));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n692_), .B2(new_n274_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT48), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n695_), .A3(new_n274_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n688_), .A2(new_n700_), .A3(new_n340_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT49), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n692_), .A2(new_n340_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G71gat), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT49), .B(new_n700_), .C1(new_n692_), .C2(new_n340_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT107), .Z(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n692_), .B2(new_n413_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT50), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n688_), .A2(new_n708_), .A3(new_n413_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1335gat));
  NOR2_X1   g511(.A1(new_n646_), .A2(new_n633_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n687_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n466_), .B1(new_n714_), .B2(new_n373_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT108), .Z(new_n716_));
  NOR3_X1   g515(.A1(new_n642_), .A2(new_n644_), .A3(KEYINPUT109), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n581_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n646_), .A2(new_n463_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n373_), .A2(new_n466_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n716_), .B1(new_n724_), .B2(new_n725_), .ZN(G1336gat));
  INV_X1    g525(.A(new_n714_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(new_n467_), .A3(new_n274_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n720_), .A2(new_n275_), .A3(new_n723_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n467_), .ZN(G1337gat));
  OAI21_X1  g529(.A(new_n722_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G99gat), .B1(new_n731_), .B2(new_n416_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n340_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n714_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT51), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n732_), .B(new_n736_), .C1(new_n714_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n487_), .A3(new_n413_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n413_), .B(new_n722_), .C1(new_n642_), .C2(new_n644_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(G106gat), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G106gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g544(.A1(new_n318_), .A2(new_n416_), .A3(new_n373_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n556_), .B(new_n530_), .C1(new_n532_), .C2(new_n540_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n551_), .B1(new_n749_), .B2(KEYINPUT112), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n550_), .A2(new_n751_), .A3(new_n530_), .A4(new_n556_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n530_), .B1(new_n532_), .B2(new_n540_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n554_), .B(new_n529_), .C1(new_n502_), .C2(new_n522_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT112), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AND4_X1   g555(.A1(new_n748_), .A2(new_n756_), .A3(new_n752_), .A4(new_n536_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n753_), .A2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n754_), .A2(new_n536_), .A3(new_n755_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT55), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n557_), .A2(KEYINPUT111), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT56), .B(new_n564_), .C1(new_n758_), .C2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n564_), .B1(new_n758_), .B2(new_n764_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n564_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n756_), .A2(new_n752_), .A3(new_n536_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT113), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n750_), .A2(new_n748_), .A3(new_n752_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n763_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n762_), .B1(new_n557_), .B2(KEYINPUT111), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n770_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n778_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n765_), .B1(new_n769_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n538_), .A2(new_n557_), .A3(new_n559_), .A4(new_n770_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n463_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n781_), .A3(new_n784_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n768_), .B(new_n770_), .C1(new_n774_), .C2(new_n777_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT114), .B1(new_n778_), .B2(KEYINPUT56), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n764_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n766_), .B(new_n768_), .C1(new_n788_), .C2(new_n770_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT115), .B1(new_n790_), .B2(new_n783_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n445_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n449_), .B(new_n792_), .C1(new_n450_), .C2(new_n452_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n459_), .C1(new_n792_), .C2(new_n444_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n565_), .A2(new_n462_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n785_), .A2(new_n791_), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT57), .A3(new_n602_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n782_), .A2(new_n462_), .A3(new_n794_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n799_), .B1(new_n801_), .B2(new_n765_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n778_), .A2(new_n800_), .A3(KEYINPUT56), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n798_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n768_), .B1(new_n788_), .B2(new_n770_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT116), .A3(new_n765_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n799_), .ZN(new_n807_));
  AND4_X1   g606(.A1(new_n798_), .A2(new_n806_), .A3(new_n803_), .A4(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n605_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n797_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT57), .B1(new_n796_), .B2(new_n602_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n581_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n684_), .A2(new_n464_), .A3(new_n567_), .A4(new_n568_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT54), .ZN(new_n814_));
  AOI211_X1 g613(.A(KEYINPUT59), .B(new_n747_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT120), .B(G113gat), .Z(new_n816_));
  NAND2_X1  g615(.A1(new_n463_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(KEYINPUT117), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n605_), .C1(new_n804_), .C2(new_n808_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n797_), .A3(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n581_), .B1(new_n822_), .B2(new_n811_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n747_), .B1(new_n823_), .B2(new_n814_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n818_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n813_), .B(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n796_), .A2(new_n602_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(new_n797_), .A3(new_n821_), .A4(new_n819_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n828_), .B1(new_n832_), .B2(new_n581_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n833_), .C2(new_n747_), .ZN(new_n834_));
  AOI211_X1 g633(.A(new_n815_), .B(new_n817_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n833_), .A2(new_n464_), .A3(new_n747_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT118), .B1(new_n836_), .B2(G113gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n824_), .A2(new_n463_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n835_), .A2(new_n842_), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n646_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n824_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n646_), .B(new_n815_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n844_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n824_), .A2(new_n849_), .A3(new_n721_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n581_), .B(new_n815_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n824_), .A2(new_n853_), .A3(new_n601_), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n643_), .B(new_n815_), .C1(new_n826_), .C2(new_n834_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n833_), .A2(new_n340_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n317_), .A2(new_n274_), .A3(new_n373_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n463_), .A3(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n569_), .A3(new_n858_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n858_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n581_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n863_), .B2(new_n643_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n602_), .A2(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n863_), .B2(new_n868_), .ZN(G1347gat));
  XNOR2_X1  g668(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n413_), .A2(new_n275_), .A3(new_n374_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n463_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873_), .B2(KEYINPUT121), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875_));
  AOI211_X1 g674(.A(new_n875_), .B(new_n872_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT123), .B(new_n870_), .C1(new_n874_), .C2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n229_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT123), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n870_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n874_), .A2(KEYINPUT123), .A3(new_n876_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n877_), .B(new_n878_), .C1(new_n881_), .C2(new_n882_), .ZN(G1348gat));
  INV_X1    g682(.A(new_n871_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n833_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n646_), .A2(new_n230_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(KEYINPUT124), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT124), .B1(new_n885_), .B2(new_n886_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G176gat), .B1(new_n889_), .B2(new_n569_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n887_), .A2(new_n888_), .A3(new_n890_), .ZN(G1349gat));
  NOR3_X1   g690(.A1(new_n833_), .A2(new_n581_), .A3(new_n884_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G183gat), .B1(new_n892_), .B2(new_n893_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n581_), .A2(new_n214_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n894_), .A2(new_n895_), .B1(new_n889_), .B2(new_n896_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n889_), .A2(new_n215_), .A3(new_n601_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n889_), .A2(new_n605_), .ZN(new_n899_));
  INV_X1    g698(.A(G190gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1351gat));
  NOR2_X1   g700(.A1(new_n275_), .A2(new_n408_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n857_), .A2(new_n463_), .A3(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g703(.A(new_n646_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n857_), .A2(new_n902_), .A3(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n906_), .B(new_n907_), .Z(G1353gat));
  NAND3_X1  g707(.A1(new_n857_), .A2(new_n721_), .A3(new_n902_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT63), .B(G211gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n909_), .B2(new_n912_), .ZN(G1354gat));
  NAND2_X1  g712(.A1(new_n857_), .A2(new_n902_), .ZN(new_n914_));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n643_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n857_), .A2(new_n601_), .A3(new_n902_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  AOI21_X1  g717(.A(G218gat), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT127), .B1(new_n914_), .B2(new_n602_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n916_), .B1(new_n919_), .B2(new_n920_), .ZN(G1355gat));
endmodule


