//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT10), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G85gat), .A3(G92gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(KEYINPUT9), .A3(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n212_), .A2(KEYINPUT64), .A3(new_n213_), .A4(new_n214_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n217_), .A2(new_n224_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT65), .ZN(new_n231_));
  INV_X1    g030(.A(new_n227_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n232_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n217_), .A4(new_n229_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT7), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(new_n220_), .A3(new_n223_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n226_), .A2(new_n248_), .A3(new_n227_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n232_), .B2(new_n225_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT8), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n255_), .A2(new_n245_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n250_), .A4(new_n249_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n238_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n209_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n238_), .A2(new_n208_), .A3(new_n259_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT34), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(KEYINPUT35), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT70), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT35), .A4(new_n264_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(KEYINPUT35), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n261_), .B(new_n267_), .C1(KEYINPUT70), .C2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G190gat), .B(G218gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G134gat), .B(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT36), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  OAI22_X1  g079(.A1(new_n273_), .A2(KEYINPUT71), .B1(KEYINPUT36), .B2(new_n276_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(KEYINPUT36), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n270_), .A2(new_n272_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n280_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT37), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n289_));
  XOR2_X1   g088(.A(G71gat), .B(G78gat), .Z(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n290_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(G8gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n296_), .B(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G127gat), .B(G155gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT16), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G183gat), .B(G211gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT17), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n304_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n296_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT73), .Z(new_n319_));
  NOR3_X1   g118(.A1(new_n287_), .A2(KEYINPUT74), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n285_), .B(KEYINPUT37), .ZN(new_n322_));
  INV_X1    g121(.A(new_n319_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n294_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n260_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n238_), .A2(new_n259_), .A3(new_n294_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G230gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT68), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n333_), .A3(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(KEYINPUT12), .A3(new_n327_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT12), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n260_), .A2(new_n337_), .A3(new_n325_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n330_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G120gat), .B(G148gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT5), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G176gat), .B(G204gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT13), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n335_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n347_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n320_), .A2(new_n324_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT18), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  AND2_X1   g155(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(G197gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT89), .B1(new_n364_), .B2(G204gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n366_));
  INV_X1    g165(.A(G204gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(G197gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(G204gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n365_), .A2(new_n368_), .A3(new_n362_), .A4(new_n369_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(new_n361_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT88), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G197gat), .B(G204gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n362_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n367_), .A2(G197gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n369_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(KEYINPUT88), .A3(KEYINPUT21), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n373_), .A2(new_n380_), .A3(KEYINPUT90), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT90), .B1(new_n373_), .B2(new_n380_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n371_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(KEYINPUT80), .A2(G183gat), .A3(G190gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n390_));
  OAI22_X1  g189(.A1(new_n388_), .A2(new_n389_), .B1(new_n390_), .B2(new_n384_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT77), .B(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(G183gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396_));
  AOI21_X1  g195(.A(G176gat), .B1(new_n396_), .B2(KEYINPUT22), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G169gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT24), .ZN(new_n400_));
  INV_X1    g199(.A(G169gat), .ZN(new_n401_));
  INV_X1    g200(.A(G176gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n401_), .A2(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n388_), .A2(new_n389_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n390_), .A2(new_n384_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n392_), .A2(KEYINPUT26), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT25), .B(G183gat), .ZN(new_n411_));
  INV_X1    g210(.A(G190gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT78), .B(KEYINPUT26), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n410_), .B(new_n411_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n399_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n383_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT94), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT94), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n383_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT26), .B(G190gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n411_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n391_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n407_), .A2(new_n408_), .B1(new_n393_), .B2(new_n412_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT22), .B(G169gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n404_), .B1(new_n425_), .B2(new_n402_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n423_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT20), .B1(new_n383_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n418_), .A2(new_n420_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n429_), .A2(new_n430_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n360_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n383_), .B2(new_n428_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n395_), .A2(new_n398_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n437_), .B(new_n371_), .C1(new_n382_), .C2(new_n381_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n434_), .B1(new_n439_), .B2(new_n359_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(KEYINPUT98), .A3(new_n360_), .A4(new_n438_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n357_), .B1(new_n433_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT99), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT99), .B(new_n357_), .C1(new_n433_), .C2(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(G155gat), .A2(G162gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(KEYINPUT1), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n448_), .A2(KEYINPUT1), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G127gat), .B(G134gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G113gat), .B(G120gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n456_), .B(KEYINPUT2), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT3), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n458_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n458_), .A2(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT3), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n449_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n448_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n460_), .A2(new_n465_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477_));
  INV_X1    g276(.A(new_n464_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n461_), .A2(new_n462_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n463_), .A2(KEYINPUT85), .A3(new_n464_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n460_), .A2(new_n474_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT4), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n460_), .A2(new_n474_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n481_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G29gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G85gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT0), .B(G57gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n475_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n484_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n498_), .B1(new_n499_), .B2(KEYINPUT100), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n501_));
  AOI211_X1 g300(.A(new_n501_), .B(new_n495_), .C1(new_n491_), .C2(new_n497_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n418_), .A2(new_n420_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n429_), .A2(new_n359_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n439_), .A2(new_n359_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(new_n357_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n356_), .A3(new_n507_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n356_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT95), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n499_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n484_), .B1(new_n496_), .B2(KEYINPUT96), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(KEYINPUT96), .B2(new_n496_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n483_), .A2(new_n490_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n518_), .B(new_n495_), .C1(new_n485_), .C2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n499_), .A2(new_n515_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n516_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n447_), .A2(new_n510_), .B1(new_n513_), .B2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n487_), .B(KEYINPUT31), .Z(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G43gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n416_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n437_), .A2(new_n528_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n211_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n399_), .A2(new_n415_), .A3(new_n528_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n528_), .B1(new_n399_), .B2(new_n415_), .ZN(new_n534_));
  OAI21_X1  g333(.A(G99gat), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G227gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(G71gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n532_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n538_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n211_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n533_), .A2(new_n534_), .A3(G99gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n532_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n527_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n541_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n543_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n526_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n486_), .A2(KEYINPUT29), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT28), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n556_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G22gat), .B(G50gat), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n383_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n474_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n459_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT29), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n383_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G228gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n383_), .B(new_n569_), .C1(new_n564_), .C2(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G78gat), .B(G106gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n573_), .A2(new_n574_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n563_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n577_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n575_), .A2(new_n582_), .A3(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n561_), .A2(new_n562_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n581_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT93), .B(new_n563_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n554_), .B(new_n580_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n523_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n580_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n554_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n580_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n578_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n582_), .B2(new_n579_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n585_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n587_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT93), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n586_), .A2(new_n581_), .A3(new_n587_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n554_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n593_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n491_), .A2(new_n497_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n495_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n501_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n499_), .A2(KEYINPUT100), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT101), .A4(new_n498_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n356_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n614_), .B1(new_n433_), .B2(new_n442_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n506_), .A2(new_n356_), .A3(new_n507_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT102), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT102), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT27), .B(new_n615_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n513_), .B2(KEYINPUT27), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n508_), .A2(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n616_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT27), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT103), .A3(new_n624_), .ZN(new_n625_));
  AND4_X1   g424(.A1(new_n613_), .A2(new_n619_), .A3(new_n621_), .A4(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n591_), .B1(new_n604_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n313_), .A2(new_n208_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n313_), .A2(new_n208_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n209_), .A2(new_n305_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT75), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT75), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n209_), .A2(new_n636_), .A3(new_n305_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n632_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n629_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n633_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G113gat), .B(G141gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G169gat), .B(G197gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n643_), .B(new_n644_), .Z(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT76), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(KEYINPUT76), .B2(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n627_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n352_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653_));
  INV_X1    g452(.A(new_n613_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n298_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n652_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n652_), .B2(new_n655_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(KEYINPUT38), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n318_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n351_), .A2(new_n650_), .A3(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT105), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n285_), .B(KEYINPUT106), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n627_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G1gat), .B1(new_n665_), .B2(new_n613_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT38), .B1(new_n656_), .B2(new_n657_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT107), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT107), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n658_), .B(new_n666_), .C1(new_n668_), .C2(new_n669_), .ZN(G1324gat));
  AND2_X1   g469(.A1(new_n621_), .A2(new_n625_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n619_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G8gat), .B1(new_n665_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n352_), .A2(new_n297_), .A3(new_n672_), .A4(new_n651_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n665_), .B2(new_n554_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT41), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n652_), .A2(G15gat), .A3(new_n554_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1326gat));
  OAI21_X1  g482(.A(G22gat), .B1(new_n665_), .B2(new_n601_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT42), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n601_), .A2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n652_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n285_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n319_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n351_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n651_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n651_), .A2(KEYINPUT110), .A3(new_n690_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n654_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n599_), .A2(new_n600_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n602_), .B1(new_n697_), .B2(new_n580_), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n594_), .B(new_n554_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n626_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n523_), .A2(new_n590_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n322_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT109), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(KEYINPUT43), .C1(new_n627_), .C2(new_n322_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n703_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n351_), .A2(new_n650_), .A3(new_n323_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n709_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(G29gat), .A3(new_n654_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n696_), .B1(new_n712_), .B2(new_n714_), .ZN(G1328gat));
  NOR2_X1   g514(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n673_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n695_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n693_), .A2(new_n694_), .A3(new_n718_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT45), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n716_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT112), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n713_), .A2(new_n672_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n708_), .B2(new_n709_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G36gat), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n722_), .A2(new_n723_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n723_), .B1(new_n722_), .B2(new_n726_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n730_));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n554_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n713_), .A2(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n733_), .B2(new_n725_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n712_), .A2(KEYINPUT113), .A3(new_n713_), .A4(new_n732_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n695_), .A2(new_n602_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n731_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT47), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT47), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n741_), .A3(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1330gat));
  AOI21_X1  g542(.A(G50gat), .B1(new_n695_), .B2(new_n592_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n713_), .A2(G50gat), .A3(new_n592_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n712_), .B2(new_n745_), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n627_), .A2(new_n649_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n349_), .A2(new_n350_), .ZN(new_n749_));
  NOR4_X1   g548(.A1(new_n748_), .A2(new_n324_), .A3(new_n749_), .A4(new_n320_), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n654_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n319_), .A2(new_n649_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n664_), .A2(new_n351_), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n613_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1332gat));
  OAI21_X1  g555(.A(G64gat), .B1(new_n754_), .B2(new_n673_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT48), .ZN(new_n758_));
  INV_X1    g557(.A(G64gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n750_), .A2(new_n759_), .A3(new_n672_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n754_), .B2(new_n554_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n750_), .A2(new_n537_), .A3(new_n602_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n754_), .B2(new_n601_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n601_), .A2(G78gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT114), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n750_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n748_), .A2(new_n749_), .A3(new_n689_), .ZN(new_n772_));
  INV_X1    g571(.A(G85gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n654_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n749_), .A2(new_n649_), .A3(new_n323_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n708_), .A2(new_n654_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n774_), .B1(new_n776_), .B2(new_n773_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT115), .ZN(G1336gat));
  INV_X1    g577(.A(G92gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n772_), .A2(new_n779_), .A3(new_n672_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n708_), .A2(new_n672_), .A3(new_n775_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n779_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT116), .ZN(G1337gat));
  NAND4_X1  g582(.A1(new_n772_), .A2(new_n602_), .A3(new_n212_), .A4(new_n214_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n708_), .A2(new_n602_), .A3(new_n775_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n211_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n772_), .A2(new_n213_), .A3(new_n592_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n708_), .A2(new_n592_), .A3(new_n775_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g593(.A1(new_n671_), .A2(new_n654_), .A3(new_n619_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n699_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT121), .B1(new_n795_), .B2(new_n603_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n628_), .A2(new_n639_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n638_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n645_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n631_), .B2(new_n639_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(KEYINPUT119), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n801_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n805_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n807_), .A2(new_n810_), .B1(new_n645_), .B2(new_n641_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n348_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n336_), .A2(new_n330_), .A3(new_n338_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n339_), .B2(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n327_), .A2(KEYINPUT12), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n294_), .B1(new_n238_), .B2(new_n259_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n338_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT55), .B(new_n329_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT118), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n329_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n820_), .A4(new_n814_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n344_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n345_), .C1(new_n822_), .C2(new_n827_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n813_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n813_), .B(KEYINPUT58), .C1(new_n829_), .C2(new_n831_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n287_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n348_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n811_), .B1(new_n348_), .B2(new_n346_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n841_), .B2(new_n285_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT57), .B(new_n688_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n836_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n836_), .B(KEYINPUT120), .C1(new_n842_), .C2(new_n843_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n659_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n749_), .A2(new_n850_), .A3(new_n753_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n323_), .A2(new_n650_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n852_), .B2(new_n351_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n849_), .B1(new_n854_), .B2(new_n322_), .ZN(new_n855_));
  AOI211_X1 g654(.A(KEYINPUT54), .B(new_n287_), .C1(new_n851_), .C2(new_n853_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n800_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n649_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n858_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT59), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n798_), .A2(KEYINPUT122), .A3(new_n799_), .ZN(new_n862_));
  AOI21_X1  g661(.A(KEYINPUT122), .B1(new_n798_), .B2(new_n799_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT59), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n855_), .A2(new_n856_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n844_), .A2(new_n319_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n862_), .B(new_n864_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n861_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n649_), .A2(G113gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT123), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n859_), .B1(new_n869_), .B2(new_n871_), .ZN(G1340gat));
  OAI21_X1  g671(.A(G120gat), .B1(new_n868_), .B2(new_n749_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n874_));
  AOI21_X1  g673(.A(G120gat), .B1(new_n351_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n874_), .B2(G120gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n858_), .A2(new_n876_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n873_), .A2(new_n879_), .ZN(G1341gat));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n318_), .B(new_n867_), .C1(new_n858_), .C2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(G127gat), .ZN(new_n883_));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n858_), .A2(new_n884_), .A3(new_n323_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT125), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(new_n888_), .A3(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1342gat));
  OAI21_X1  g689(.A(G134gat), .B1(new_n868_), .B2(new_n322_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n662_), .A2(G134gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n860_), .B2(new_n892_), .ZN(G1343gat));
  AOI21_X1  g692(.A(new_n593_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(KEYINPUT126), .A3(new_n796_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT126), .B1(new_n894_), .B2(new_n796_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n649_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G141gat), .ZN(new_n899_));
  INV_X1    g698(.A(G141gat), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(new_n649_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1344gat));
  OAI21_X1  g701(.A(new_n351_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G148gat), .ZN(new_n904_));
  INV_X1    g703(.A(G148gat), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n351_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1345gat));
  OAI21_X1  g706(.A(new_n323_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n323_), .B(new_n911_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1346gat));
  INV_X1    g712(.A(G162gat), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n914_), .B(new_n663_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n897_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n322_), .B1(new_n916_), .B2(new_n895_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n917_), .B2(new_n914_), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n866_), .A2(new_n865_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n673_), .A2(new_n654_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n602_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n601_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n919_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925_), .B2(new_n650_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n924_), .A2(new_n649_), .A3(new_n425_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n927_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n924_), .B2(new_n351_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n592_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n921_), .A2(new_n402_), .A3(new_n749_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1349gat));
  NOR3_X1   g734(.A1(new_n925_), .A2(new_n411_), .A3(new_n659_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n323_), .A3(new_n922_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n393_), .B2(new_n937_), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n925_), .B2(new_n322_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n924_), .A2(new_n421_), .A3(new_n663_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n848_), .A2(new_n857_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n698_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n920_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n649_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n351_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g748(.A1(new_n943_), .A2(new_n659_), .A3(new_n944_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n953_), .B1(new_n950_), .B2(new_n951_), .ZN(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n894_), .A2(new_n955_), .A3(new_n663_), .A4(new_n920_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n943_), .A2(new_n322_), .A3(new_n944_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n957_), .B2(new_n955_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  OAI211_X1 g759(.A(KEYINPUT127), .B(new_n956_), .C1(new_n957_), .C2(new_n955_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1355gat));
endmodule


