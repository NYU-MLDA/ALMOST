//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n970_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_;
  INV_X1    g000(.A(KEYINPUT8), .ZN(new_n202_));
  AND2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR3_X1   g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n203_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT66), .B1(new_n217_), .B2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n214_), .A2(new_n215_), .A3(new_n203_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n203_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n209_), .A2(new_n216_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n202_), .A2(new_n224_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  INV_X1    g041(.A(G99gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n226_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n210_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n232_), .A2(new_n233_), .A3(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n241_), .B1(new_n246_), .B2(new_n222_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n217_), .A2(KEYINPUT66), .A3(new_n223_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(KEYINPUT8), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G78gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT11), .ZN(new_n252_));
  XOR2_X1   g051(.A(G71gat), .B(G78gat), .Z(new_n253_));
  INV_X1    g052(.A(G64gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G57gat), .ZN(new_n255_));
  INV_X1    g054(.A(G57gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G64gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n257_), .A3(KEYINPUT11), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n252_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n240_), .A2(new_n249_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT67), .B(new_n252_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(KEYINPUT12), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n266_), .B1(new_n240_), .B2(new_n249_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n217_), .A2(KEYINPUT66), .A3(new_n223_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n270_), .A2(new_n224_), .A3(new_n202_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n236_), .A2(new_n239_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n241_), .B(new_n202_), .C1(new_n246_), .C2(new_n222_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n269_), .B1(new_n275_), .B2(new_n261_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G230gat), .A2(G233gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n261_), .B1(new_n240_), .B2(new_n249_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n262_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G120gat), .B(G148gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT5), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G176gat), .B(G204gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n264_), .A2(KEYINPUT12), .A3(new_n265_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n240_), .A2(new_n249_), .A3(new_n261_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n290_), .B(new_n291_), .C1(new_n280_), .C2(KEYINPUT12), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n281_), .B(new_n288_), .C1(new_n292_), .C2(new_n279_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n295_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n287_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(new_n294_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT69), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(new_n282_), .A3(new_n286_), .A4(new_n296_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n299_), .A2(new_n302_), .A3(KEYINPUT13), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT13), .B1(new_n299_), .B2(new_n302_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT70), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307_));
  XOR2_X1   g106(.A(G29gat), .B(G36gat), .Z(new_n308_));
  XOR2_X1   g107(.A(G43gat), .B(G50gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G29gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G43gat), .B(G50gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(KEYINPUT75), .A3(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G1gat), .B(G8gat), .Z(new_n319_));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G1gat), .B(G8gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT72), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G15gat), .B(G22gat), .ZN(new_n325_));
  INV_X1    g124(.A(G1gat), .ZN(new_n326_));
  INV_X1    g125(.A(G8gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT14), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n321_), .A3(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n318_), .A2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n316_), .A2(new_n330_), .A3(new_n317_), .A4(new_n332_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT76), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G229gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n318_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n314_), .B(KEYINPUT15), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n333_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n337_), .A3(new_n335_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G169gat), .B(G197gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  AND3_X1   g146(.A1(new_n341_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n307_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(new_n344_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n347_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n341_), .A2(new_n344_), .A3(new_n347_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(KEYINPUT77), .A3(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n303_), .A2(new_n304_), .A3(KEYINPUT70), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n306_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT22), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  OR3_X1    g162(.A1(new_n360_), .A2(KEYINPUT80), .A3(KEYINPUT22), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT81), .B(G176gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT80), .B1(new_n360_), .B2(KEYINPUT22), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT78), .B(G190gat), .Z(new_n368_));
  INV_X1    g167(.A(G183gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT23), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n370_), .A2(new_n372_), .B1(G169gat), .B2(G176gat), .ZN(new_n373_));
  INV_X1    g172(.A(G176gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n360_), .A2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT24), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(KEYINPUT24), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n368_), .A2(KEYINPUT26), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT25), .B(G183gat), .ZN(new_n382_));
  INV_X1    g181(.A(G190gat), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT26), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n367_), .A2(new_n373_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT88), .ZN(new_n388_));
  INV_X1    g187(.A(G197gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G204gat), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n388_), .B(KEYINPUT21), .C1(KEYINPUT88), .C2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G211gat), .B(G218gat), .Z(new_n392_));
  INV_X1    g191(.A(KEYINPUT21), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n387_), .ZN(new_n394_));
  INV_X1    g193(.A(G204gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G197gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT21), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT89), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n392_), .A2(new_n401_), .A3(KEYINPUT21), .A4(new_n397_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n391_), .A2(new_n394_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n359_), .B1(new_n386_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n383_), .A2(KEYINPUT26), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n382_), .A2(new_n384_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n380_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT92), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n372_), .B1(G183gat), .B2(G190gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n377_), .B(KEYINPUT93), .Z(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT22), .B(G169gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n365_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n411_), .A2(KEYINPUT94), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT94), .B1(new_n411_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n410_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n380_), .A2(KEYINPUT92), .A3(new_n406_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n391_), .A2(new_n394_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n400_), .A2(new_n402_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n404_), .A2(KEYINPUT91), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT19), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n373_), .A2(new_n367_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n380_), .A2(new_n385_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT20), .B1(new_n428_), .B2(new_n421_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n421_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n416_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n424_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G8gat), .B(G36gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT18), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G64gat), .B(G92gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n440_), .B(new_n441_), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n404_), .A2(KEYINPUT91), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n418_), .A2(new_n421_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n431_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n424_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n409_), .A2(new_n416_), .A3(new_n403_), .A4(new_n417_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(new_n433_), .A3(KEYINPUT20), .A4(new_n425_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n442_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(KEYINPUT27), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT102), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT102), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n444_), .A2(new_n451_), .A3(new_n454_), .A4(KEYINPUT27), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G155gat), .A2(G162gat), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n457_), .A2(KEYINPUT1), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n459_), .B2(KEYINPUT1), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n461_), .B2(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G141gat), .A2(G148gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n467_), .B(KEYINPUT3), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n472_), .B(new_n473_), .C1(KEYINPUT2), .C2(new_n466_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G155gat), .B(G162gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT86), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT29), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(G228gat), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n479_), .A2(new_n421_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n469_), .B2(new_n477_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n487_), .B2(new_n403_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G78gat), .B(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n484_), .A2(new_n488_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n469_), .A2(new_n477_), .A3(new_n486_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n463_), .A2(new_n468_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT28), .B1(new_n497_), .B2(new_n486_), .ZN(new_n498_));
  OAI21_X1  g297(.A(G22gat), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n495_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(KEYINPUT28), .A3(new_n486_), .ZN(new_n501_));
  INV_X1    g300(.A(G22gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(G50gat), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n493_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(G50gat), .B1(new_n499_), .B2(new_n503_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n491_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n490_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n505_), .A2(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n499_), .A2(new_n503_), .ZN(new_n511_));
  INV_X1    g310(.A(G50gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n510_), .A2(new_n513_), .A3(new_n493_), .A4(new_n504_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n448_), .A2(KEYINPUT95), .A3(new_n442_), .A4(new_n450_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n425_), .B1(new_n422_), .B2(new_n431_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n450_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n443_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n447_), .B2(new_n424_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT95), .B1(new_n522_), .B2(new_n442_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n516_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n456_), .A2(new_n515_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G120gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G127gat), .B(G134gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n528_), .A2(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n527_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G134gat), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT82), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n530_), .A3(new_n526_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n478_), .B2(KEYINPUT96), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n531_), .A2(new_n532_), .A3(new_n527_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n526_), .B1(new_n535_), .B2(new_n530_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n497_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(KEYINPUT4), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n497_), .B2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n478_), .A2(KEYINPUT97), .A3(new_n546_), .A4(new_n537_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G225gat), .A2(G233gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n544_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT98), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT98), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n544_), .A2(new_n550_), .A3(new_n555_), .A4(new_n552_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n538_), .A2(new_n543_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n551_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n554_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G1gat), .B(G29gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G85gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n554_), .A2(new_n566_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G71gat), .B(G99gat), .ZN(new_n569_));
  INV_X1    g368(.A(G43gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n386_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n537_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G227gat), .A2(G233gat), .ZN(new_n574_));
  INV_X1    g373(.A(G15gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT30), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT31), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n573_), .B(new_n578_), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n568_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n525_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT103), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n565_), .A2(new_n567_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n515_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n456_), .A2(new_n582_), .A3(new_n524_), .A4(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n524_), .A2(new_n453_), .A3(new_n455_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n515_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n568_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT103), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n442_), .A2(KEYINPUT32), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n432_), .B2(new_n437_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n522_), .B2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n567_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n451_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n538_), .A2(new_n543_), .A3(new_n552_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n564_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT100), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n544_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(KEYINPUT100), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n597_), .A2(new_n603_), .A3(new_n520_), .A4(new_n517_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n593_), .B1(new_n595_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n515_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n585_), .A2(new_n589_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n579_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n581_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n358_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n240_), .A2(new_n249_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n342_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n314_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n612_), .B(new_n617_), .C1(new_n618_), .C2(new_n611_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n615_), .A2(new_n616_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT71), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n611_), .B2(new_n618_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n619_), .B(new_n620_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n342_), .B2(new_n611_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n622_), .B2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(KEYINPUT36), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n623_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n629_), .B(KEYINPUT36), .Z(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT37), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n623_), .A2(new_n626_), .A3(new_n630_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n623_), .A2(new_n626_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n636_), .B(new_n637_), .C1(new_n638_), .C2(new_n633_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n333_), .B(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT73), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n264_), .A2(new_n265_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(G127gat), .B(G155gat), .Z(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G183gat), .B(G211gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n643_), .A2(new_n644_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n645_), .A2(KEYINPUT17), .A3(new_n651_), .A4(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n642_), .A2(new_n261_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n642_), .A2(new_n261_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n650_), .B(KEYINPUT17), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n654_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n640_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n610_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n326_), .A3(new_n583_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n306_), .A2(new_n357_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n658_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(KEYINPUT104), .A3(new_n356_), .A4(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n637_), .B1(new_n638_), .B2(new_n633_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n609_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n672_), .B1(new_n358_), .B2(new_n658_), .ZN(new_n673_));
  AND4_X1   g472(.A1(new_n583_), .A2(new_n668_), .A3(new_n671_), .A4(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n663_), .B(new_n664_), .C1(new_n326_), .C2(new_n674_), .ZN(G1324gat));
  NAND4_X1  g474(.A1(new_n668_), .A2(new_n586_), .A3(new_n673_), .A4(new_n671_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G8gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n610_), .A2(new_n327_), .A3(new_n586_), .A4(new_n659_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT105), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n679_), .A2(new_n681_), .A3(KEYINPUT40), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  NAND3_X1  g486(.A1(new_n660_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n668_), .A2(new_n579_), .A3(new_n673_), .A4(new_n671_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT41), .B1(new_n689_), .B2(G15gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(G1326gat));
  NAND3_X1  g491(.A1(new_n660_), .A2(new_n502_), .A3(new_n587_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n668_), .A2(new_n587_), .A3(new_n673_), .A4(new_n671_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(G22gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n694_), .B2(G22gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1327gat));
  NOR2_X1   g497(.A1(new_n667_), .A2(new_n669_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n610_), .A2(new_n699_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n700_), .A2(G29gat), .A3(new_n568_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n635_), .A2(new_n639_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n702_), .B2(KEYINPUT106), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n704_), .B1(new_n609_), .B2(new_n702_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n584_), .A2(new_n524_), .A3(new_n455_), .A4(new_n453_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n706_), .A2(KEYINPUT103), .B1(new_n605_), .B2(new_n515_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n579_), .B1(new_n707_), .B2(new_n585_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n640_), .B(new_n703_), .C1(new_n708_), .C2(new_n581_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n306_), .A2(new_n356_), .A3(new_n357_), .A4(new_n658_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n714_), .B(new_n711_), .C1(new_n705_), .C2(new_n709_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n713_), .A2(new_n715_), .A3(new_n568_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G29gat), .B1(new_n716_), .B2(new_n717_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n701_), .B1(new_n718_), .B2(new_n719_), .ZN(G1328gat));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  INV_X1    g520(.A(G36gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n713_), .A2(new_n715_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n586_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n610_), .A2(new_n722_), .A3(new_n586_), .A4(new_n699_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT45), .Z(new_n726_));
  OAI21_X1  g525(.A(new_n721_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n725_), .B(KEYINPUT45), .ZN(new_n728_));
  INV_X1    g527(.A(new_n586_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n713_), .A2(new_n715_), .A3(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n728_), .B(KEYINPUT46), .C1(new_n730_), .C2(new_n722_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(G1329gat));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n570_), .B1(new_n723_), .B2(new_n579_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n700_), .A2(G43gat), .A3(new_n608_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n735_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n713_), .A2(new_n715_), .A3(new_n608_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT47), .B(new_n737_), .C1(new_n738_), .C2(new_n570_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1330gat));
  INV_X1    g539(.A(new_n700_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G50gat), .B1(new_n741_), .B2(new_n587_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n515_), .A2(new_n512_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n723_), .B2(new_n743_), .ZN(G1331gat));
  INV_X1    g543(.A(new_n609_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n356_), .B1(new_n306_), .B2(new_n357_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n659_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n568_), .B1(new_n749_), .B2(KEYINPUT108), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(KEYINPUT108), .B2(new_n749_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n671_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n356_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n665_), .A2(new_n753_), .A3(new_n667_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n752_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n568_), .A2(new_n256_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n751_), .A2(new_n256_), .B1(new_n758_), .B2(new_n759_), .ZN(G1332gat));
  NAND3_X1  g559(.A1(new_n749_), .A2(new_n254_), .A3(new_n586_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n586_), .A3(new_n757_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G64gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G64gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1333gat));
  OR3_X1    g565(.A1(new_n748_), .A2(G71gat), .A3(new_n608_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n579_), .A3(new_n757_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G71gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G71gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1334gat));
  OR3_X1    g571(.A1(new_n748_), .A2(G78gat), .A3(new_n515_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n756_), .A2(new_n587_), .A3(new_n757_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G78gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n746_), .A2(new_n658_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n710_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n568_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n747_), .A2(new_n699_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n583_), .A2(new_n218_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(G1336gat));
  OAI21_X1  g584(.A(G92gat), .B1(new_n781_), .B2(new_n729_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n586_), .A2(new_n219_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n783_), .B2(new_n787_), .ZN(G1337gat));
  AOI21_X1  g587(.A(new_n779_), .B1(new_n709_), .B2(new_n705_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n243_), .B1(new_n789_), .B2(new_n579_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n579_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n783_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1338gat));
  NOR2_X1   g594(.A1(new_n781_), .A2(new_n515_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n226_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n515_), .A2(G106gat), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n745_), .A2(new_n746_), .A3(new_n699_), .A4(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n226_), .B1(new_n789_), .B2(new_n587_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(KEYINPUT52), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT53), .B1(new_n798_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n797_), .B1(new_n796_), .B2(new_n226_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(KEYINPUT52), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .A4(new_n802_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n805_), .A2(new_n809_), .ZN(G1339gat));
  NAND4_X1  g609(.A1(new_n729_), .A2(new_n583_), .A3(new_n515_), .A4(new_n579_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT116), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT111), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n292_), .B2(new_n279_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n292_), .A2(new_n279_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n292_), .A2(new_n817_), .A3(new_n279_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n286_), .B(new_n816_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n350_), .A2(new_n355_), .A3(new_n293_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n277_), .B1(new_n268_), .B2(new_n276_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n278_), .B1(new_n825_), .B2(new_n817_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n821_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n816_), .B1(new_n828_), .B2(new_n286_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n813_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n286_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n815_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(KEYINPUT112), .A3(new_n822_), .A4(new_n823_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n335_), .A2(new_n338_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n347_), .B1(new_n835_), .B2(new_n343_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n336_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n834_), .B1(new_n354_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n354_), .A2(new_n838_), .A3(new_n834_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n299_), .A2(new_n302_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n830_), .A2(new_n833_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n669_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(KEYINPUT57), .A3(new_n669_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n841_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n293_), .B1(new_n852_), .B2(new_n839_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n288_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n814_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n831_), .A2(KEYINPUT56), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n851_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n849_), .B1(new_n857_), .B2(new_n702_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n293_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n831_), .B2(KEYINPUT56), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n854_), .A2(new_n814_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n850_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(KEYINPUT115), .A3(new_n640_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n855_), .A2(KEYINPUT58), .A3(new_n856_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n858_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n847_), .A2(new_n848_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n658_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n356_), .B(new_n658_), .C1(new_n635_), .C2(new_n639_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n305_), .B2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n870_), .B(new_n869_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n871_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n812_), .B1(new_n868_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT117), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n871_), .A2(new_n873_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n658_), .B2(new_n867_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n878_), .B(KEYINPUT59), .C1(new_n880_), .C2(new_n812_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n867_), .A2(KEYINPUT118), .A3(new_n658_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n874_), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT118), .B1(new_n867_), .B2(new_n658_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT119), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n883_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n882_), .A2(new_n888_), .A3(new_n356_), .A4(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G113gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n875_), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n893_), .A2(G113gat), .A3(new_n753_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1340gat));
  NAND4_X1  g694(.A1(new_n882_), .A2(new_n888_), .A3(new_n665_), .A4(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G120gat), .ZN(new_n897_));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n666_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n875_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(G1341gat));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n658_), .A2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT120), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n882_), .A2(new_n888_), .A3(new_n890_), .A4(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n893_), .B2(new_n658_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1342gat));
  NAND4_X1  g706(.A1(new_n882_), .A2(new_n888_), .A3(new_n640_), .A4(new_n890_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G134gat), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n893_), .A2(G134gat), .A3(new_n669_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1343gat));
  NAND2_X1  g710(.A1(new_n868_), .A2(new_n874_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n579_), .A2(new_n515_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n586_), .A2(new_n568_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n753_), .ZN(new_n917_));
  INV_X1    g716(.A(G141gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1344gat));
  NOR2_X1   g718(.A1(new_n916_), .A2(new_n666_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT121), .B(G148gat), .Z(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1345gat));
  NOR2_X1   g721(.A1(new_n916_), .A2(new_n658_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT61), .B(G155gat), .Z(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  AND2_X1   g724(.A1(new_n914_), .A2(new_n915_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G162gat), .B1(new_n926_), .B2(new_n670_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n640_), .A2(G162gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT122), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n926_), .B2(new_n929_), .ZN(G1347gat));
  OR2_X1    g729(.A1(new_n885_), .A2(new_n886_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n729_), .A2(new_n580_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n587_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n931_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n356_), .A2(new_n412_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT124), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n356_), .B(new_n934_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n360_), .B1(new_n940_), .B2(KEYINPUT62), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n939_), .B(new_n941_), .C1(new_n940_), .C2(KEYINPUT62), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n939_), .A2(new_n941_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n943_), .A2(KEYINPUT123), .A3(new_n944_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n938_), .A2(new_n942_), .A3(new_n945_), .ZN(G1348gat));
  NAND2_X1  g745(.A1(new_n935_), .A2(new_n665_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n880_), .A2(new_n587_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n666_), .A2(new_n374_), .A3(new_n933_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n947_), .A2(new_n365_), .B1(new_n948_), .B2(new_n949_), .ZN(G1349gat));
  NOR2_X1   g749(.A1(new_n658_), .A2(new_n382_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n948_), .A2(new_n667_), .A3(new_n932_), .ZN(new_n952_));
  AOI22_X1  g751(.A1(new_n935_), .A2(new_n951_), .B1(new_n369_), .B2(new_n952_), .ZN(G1350gat));
  NAND4_X1  g752(.A1(new_n935_), .A2(new_n384_), .A3(new_n405_), .A4(new_n670_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n931_), .A2(new_n640_), .A3(new_n934_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n955_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n954_), .B1(new_n383_), .B2(new_n956_), .ZN(G1351gat));
  NOR2_X1   g756(.A1(new_n729_), .A2(new_n583_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n912_), .A2(new_n356_), .A3(new_n913_), .A4(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n389_), .B1(new_n959_), .B2(KEYINPUT125), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n959_), .B2(KEYINPUT125), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n959_), .A2(KEYINPUT125), .A3(new_n962_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n961_), .A2(new_n964_), .A3(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n965_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n960_), .B1(new_n967_), .B2(new_n963_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1352gat));
  NAND2_X1  g768(.A1(new_n914_), .A2(new_n958_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n970_), .A2(new_n666_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(new_n395_), .ZN(G1353gat));
  AOI21_X1  g771(.A(new_n658_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  NAND4_X1  g772(.A1(new_n912_), .A2(new_n913_), .A3(new_n958_), .A4(new_n973_), .ZN(new_n974_));
  OR2_X1    g773(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n975_));
  NOR2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n977_));
  AND3_X1   g776(.A1(new_n975_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n976_), .B1(new_n975_), .B2(new_n977_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n978_), .A2(new_n979_), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n970_), .B2(new_n702_), .ZN(new_n981_));
  OR2_X1    g780(.A1(new_n669_), .A2(G218gat), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n970_), .B2(new_n982_), .ZN(G1355gat));
endmodule


