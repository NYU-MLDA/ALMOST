//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_;
  NOR2_X1   g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT89), .ZN(new_n203_));
  OR2_X1    g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n202_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n204_), .A2(new_n206_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT28), .B1(new_n220_), .B2(KEYINPUT29), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n209_), .A2(new_n208_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n202_), .A2(KEYINPUT89), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n202_), .A2(KEYINPUT89), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n225_), .A2(new_n207_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G22gat), .B(G50gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n221_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n221_), .B2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT93), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n230_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n220_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n227_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT93), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n221_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n220_), .A2(KEYINPUT29), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G211gat), .B(G218gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT92), .ZN(new_n245_));
  INV_X1    g044(.A(G204gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(G197gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(G197gat), .ZN(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(G204gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n243_), .B1(new_n253_), .B2(new_n248_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n247_), .A2(new_n250_), .A3(new_n243_), .A4(new_n248_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n242_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n252_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT90), .Z(new_n261_));
  AND3_X1   g060(.A1(new_n241_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n241_), .B2(new_n259_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n233_), .A2(new_n240_), .A3(new_n264_), .ZN(new_n265_));
  OAI221_X1 g064(.A(KEYINPUT93), .B1(new_n262_), .B2(new_n263_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G78gat), .B(G106gat), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n268_), .A3(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(G15gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT30), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278_));
  INV_X1    g077(.A(G183gat), .ZN(new_n279_));
  INV_X1    g078(.A(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n280_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT85), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n281_), .A2(KEYINPUT86), .A3(new_n282_), .A4(new_n283_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT22), .B(G169gat), .ZN(new_n291_));
  INV_X1    g090(.A(G176gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n286_), .A2(new_n289_), .A3(new_n290_), .A4(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G190gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n279_), .A2(KEYINPUT25), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(KEYINPUT83), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT25), .B(G183gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(KEYINPUT83), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G183gat), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n303_), .A2(KEYINPUT83), .A3(KEYINPUT84), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n296_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n289_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(new_n292_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n281_), .A2(new_n282_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n294_), .B1(new_n306_), .B2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G71gat), .B(G99gat), .Z(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT87), .B(G43gat), .Z(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  NOR2_X1   g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n318_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n277_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n277_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n319_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT88), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n323_), .B2(new_n319_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n320_), .A2(new_n277_), .A3(new_n321_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G127gat), .B(G134gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(G113gat), .B(G120gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT31), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  OAI211_X1 g135(.A(KEYINPUT88), .B(new_n336_), .C1(new_n322_), .C2(new_n325_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT98), .B1(new_n220_), .B2(new_n333_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n220_), .A2(new_n333_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n348_), .A2(KEYINPUT4), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n346_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n345_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n344_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT33), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT33), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n351_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n349_), .A2(new_n345_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n343_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n356_), .B1(new_n361_), .B2(new_n355_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT97), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n244_), .A2(new_n251_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n253_), .A2(new_n248_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n255_), .B1(new_n365_), .B2(new_n243_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n254_), .A2(KEYINPUT91), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n258_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n364_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n281_), .A2(new_n282_), .A3(new_n312_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n289_), .B2(new_n308_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n298_), .A2(new_n303_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n304_), .B1(new_n375_), .B2(new_n299_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n372_), .B1(new_n376_), .B2(new_n296_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n377_), .A3(new_n294_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n308_), .A2(new_n287_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n296_), .B2(new_n373_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT96), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n281_), .A2(new_n312_), .A3(new_n381_), .A4(new_n282_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(KEYINPUT96), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n293_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n258_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n386_));
  OAI22_X1  g185(.A1(new_n384_), .A2(new_n385_), .B1(new_n386_), .B2(new_n364_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n378_), .A2(new_n387_), .A3(KEYINPUT20), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n389_));
  AND2_X1   g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT95), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n363_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n315_), .B2(new_n259_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n380_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n383_), .A2(new_n382_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n385_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(new_n370_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n363_), .B(new_n392_), .C1(new_n395_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n401_), .B1(new_n398_), .B2(new_n370_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n315_), .A2(new_n259_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n391_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n394_), .A2(new_n411_), .A3(new_n400_), .A4(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n362_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n355_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n353_), .A2(new_n344_), .A3(new_n354_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n405_), .B2(KEYINPUT100), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n402_), .A2(new_n403_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n419_), .A2(new_n391_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n417_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT100), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n405_), .B2(new_n422_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n415_), .A2(new_n416_), .B1(new_n418_), .B2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n273_), .B(new_n338_), .C1(new_n414_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n400_), .A2(new_n404_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(new_n393_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n428_), .A2(new_n411_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n427_), .A2(new_n409_), .A3(new_n393_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n426_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n270_), .A2(new_n271_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n395_), .A2(new_n399_), .A3(new_n392_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n391_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n409_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT27), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT101), .B1(new_n430_), .B2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n426_), .B1(new_n420_), .B2(new_n409_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT101), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n412_), .A3(new_n439_), .ZN(new_n440_));
  AND4_X1   g239(.A1(new_n431_), .A2(new_n432_), .A3(new_n437_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n440_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT27), .B1(new_n410_), .B2(new_n412_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT102), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT102), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n431_), .A2(new_n445_), .A3(new_n437_), .A4(new_n440_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n272_), .A2(new_n338_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n441_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n415_), .A2(new_n416_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n425_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G57gat), .B(G64gat), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n452_), .A2(KEYINPUT11), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G71gat), .B(G78gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(KEYINPUT11), .B2(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n454_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G85gat), .B(G92gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT7), .ZN(new_n462_));
  NOR2_X1   g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT65), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT6), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  AOI211_X1 g273(.A(KEYINPUT8), .B(new_n460_), .C1(new_n469_), .C2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(KEYINPUT66), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n462_), .A2(new_n467_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n463_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n471_), .A2(new_n473_), .A3(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n464_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n460_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(KEYINPUT67), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT67), .B1(new_n483_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n476_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n460_), .A2(KEYINPUT9), .ZN(new_n490_));
  INV_X1    g289(.A(G92gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n460_), .B1(KEYINPUT9), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT64), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT10), .B(G99gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n474_), .B1(new_n496_), .B2(G106gat), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n488_), .A2(new_n489_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n489_), .B1(new_n488_), .B2(new_n499_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n459_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n471_), .A2(new_n473_), .A3(new_n481_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n481_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n460_), .B1(new_n506_), .B2(new_n469_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n507_), .B2(KEYINPUT67), .ZN(new_n508_));
  INV_X1    g307(.A(new_n487_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n475_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT68), .B1(new_n510_), .B2(new_n498_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n488_), .A2(new_n489_), .A3(new_n499_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n458_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n502_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G230gat), .ZN(new_n515_));
  INV_X1    g314(.A(G233gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n488_), .A2(new_n499_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(KEYINPUT12), .A3(new_n459_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n458_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n513_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n518_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G120gat), .B(G148gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n518_), .B(new_n530_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n533_), .A2(new_n535_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n536_));
  AND2_X1   g335(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n537_));
  NOR2_X1   g336(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n532_), .B(new_n534_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT81), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT78), .B(G15gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G22gat), .ZN(new_n546_));
  INV_X1    g345(.A(G1gat), .ZN(new_n547_));
  INV_X1    g346(.A(G8gat), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G1gat), .B(G8gat), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G29gat), .B(G36gat), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT73), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n556_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G43gat), .B(G50gat), .Z(new_n559_));
  OR3_X1    g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n559_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n554_), .A2(KEYINPUT80), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT80), .B1(new_n554_), .B2(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n562_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n554_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n565_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n554_), .A2(new_n562_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n566_), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n544_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n544_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n563_), .A2(new_n564_), .B1(new_n562_), .B2(new_n554_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n574_), .B(new_n575_), .C1(new_n566_), .C2(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n573_), .A2(KEYINPUT82), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT82), .B1(new_n573_), .B2(new_n577_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n451_), .A2(new_n540_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT34), .Z(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n500_), .A2(new_n501_), .A3(new_n562_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n519_), .A2(new_n568_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n584_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT74), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(KEYINPUT75), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n585_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n587_), .A2(new_n590_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n585_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n511_), .A2(new_n512_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(KEYINPUT36), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n592_), .A2(new_n596_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT76), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n592_), .A2(new_n596_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n599_), .B(KEYINPUT36), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n592_), .A2(new_n596_), .A3(KEYINPUT76), .A4(new_n600_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(KEYINPUT37), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT37), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n611_), .A3(new_n601_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n609_), .B1(new_n608_), .B2(KEYINPUT37), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n554_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n459_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G127gat), .B(G155gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT17), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT79), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT79), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n618_), .A2(new_n627_), .A3(new_n624_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n618_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n622_), .B(KEYINPUT17), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n626_), .A2(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n615_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n581_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n450_), .B(KEYINPUT103), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n547_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT38), .ZN(new_n637_));
  INV_X1    g436(.A(new_n540_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n573_), .A2(new_n577_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n606_), .A2(new_n642_), .A3(new_n601_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n606_), .B2(new_n601_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n641_), .A2(new_n451_), .A3(new_n646_), .A4(new_n631_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n450_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n637_), .A2(new_n649_), .ZN(G1324gat));
  INV_X1    g449(.A(new_n447_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n634_), .A2(new_n548_), .A3(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G8gat), .B1(new_n647_), .B2(new_n447_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n653_), .A2(KEYINPUT105), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(KEYINPUT105), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n654_), .A2(new_n655_), .A3(KEYINPUT39), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n652_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT40), .B(new_n652_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647_), .B2(new_n338_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n338_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n634_), .A2(new_n275_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(G22gat), .B1(new_n647_), .B2(new_n273_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n634_), .A2(new_n673_), .A3(new_n272_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1327gat));
  NOR2_X1   g474(.A1(new_n646_), .A2(new_n631_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n581_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(G29gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n450_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n608_), .A2(KEYINPUT37), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT77), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n684_), .A2(KEYINPUT107), .A3(new_n610_), .A4(new_n612_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n451_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n451_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(KEYINPUT44), .A3(new_n632_), .A4(new_n641_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n686_), .A2(KEYINPUT43), .B1(new_n451_), .B2(new_n689_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n641_), .A2(new_n632_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n692_), .A2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(new_n635_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n680_), .B1(new_n698_), .B2(new_n679_), .ZN(G1328gat));
  OR2_X1    g498(.A1(new_n651_), .A2(KEYINPUT109), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n651_), .A2(KEYINPUT109), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n677_), .A2(G36gat), .A3(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT45), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n692_), .A2(new_n651_), .A3(new_n696_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G36gat), .B1(new_n705_), .B2(new_n706_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT46), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1329gat));
  NOR3_X1   g512(.A1(new_n677_), .A2(G43gat), .A3(new_n338_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n692_), .A2(new_n668_), .A3(new_n696_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G43gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g516(.A(G50gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n678_), .A2(new_n718_), .A3(new_n272_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n697_), .A2(new_n272_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G50gat), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT110), .B(new_n718_), .C1(new_n697_), .C2(new_n272_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1331gat));
  INV_X1    g523(.A(new_n451_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n725_), .A2(new_n540_), .A3(new_n639_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n633_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n728_), .A2(KEYINPUT111), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(KEYINPUT111), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n635_), .A3(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n631_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n733_));
  NOR4_X1   g532(.A1(new_n725_), .A2(new_n645_), .A3(new_n540_), .A4(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n648_), .A2(new_n732_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n731_), .A2(new_n732_), .B1(new_n734_), .B2(new_n735_), .ZN(G1332gat));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  INV_X1    g536(.A(new_n702_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT48), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n728_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n734_), .B2(new_n668_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT49), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n728_), .A2(new_n743_), .A3(new_n668_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n734_), .B2(new_n272_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT50), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n728_), .A2(new_n748_), .A3(new_n272_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1335gat));
  AND2_X1   g551(.A1(new_n726_), .A2(new_n676_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n635_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT112), .Z(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n687_), .A2(new_n757_), .A3(new_n690_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n638_), .A2(new_n632_), .A3(new_n640_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n694_), .A2(new_n757_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n691_), .A2(KEYINPUT113), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(KEYINPUT114), .A3(new_n758_), .A4(new_n760_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n763_), .A2(new_n765_), .A3(G85gat), .A4(new_n450_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n755_), .A2(new_n766_), .ZN(G1336gat));
  NAND3_X1  g566(.A1(new_n753_), .A2(new_n491_), .A3(new_n651_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n763_), .A2(new_n738_), .A3(new_n765_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n491_), .ZN(G1337gat));
  NAND3_X1  g569(.A1(new_n763_), .A2(new_n668_), .A3(new_n765_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G99gat), .ZN(new_n772_));
  INV_X1    g571(.A(new_n496_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n753_), .A2(new_n668_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n772_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  INV_X1    g578(.A(G106gat), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n759_), .A2(new_n273_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n691_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n753_), .A2(new_n780_), .A3(new_n272_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g586(.A(new_n635_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n447_), .A2(new_n448_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n513_), .B(new_n520_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n517_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n500_), .A2(new_n501_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n517_), .B1(new_n797_), .B2(new_n458_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n522_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n502_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n798_), .A2(new_n800_), .A3(KEYINPUT55), .A4(new_n520_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n796_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n531_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT115), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n802_), .A2(KEYINPUT115), .A3(new_n804_), .A4(new_n531_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n639_), .A2(new_n534_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n543_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n576_), .A2(new_n566_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n566_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n574_), .B(new_n543_), .C1(new_n566_), .C2(new_n576_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n645_), .B1(new_n810_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n792_), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n802_), .A2(new_n804_), .A3(new_n531_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n535_), .A2(new_n816_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n615_), .A2(new_n825_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n808_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n817_), .B1(new_n831_), .B2(new_n807_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT116), .B(new_n830_), .C1(new_n832_), .C2(new_n645_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n820_), .A2(new_n821_), .A3(new_n829_), .A4(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n632_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n733_), .B1(new_n536_), .B2(new_n539_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n688_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n688_), .B2(new_n836_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n791_), .B1(new_n835_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n639_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n839_), .A2(new_n840_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n834_), .B2(new_n632_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n791_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n830_), .B1(new_n832_), .B2(new_n645_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n829_), .A2(new_n821_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n632_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n841_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n791_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n846_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT117), .B(G113gat), .Z(new_n855_));
  NAND2_X1  g654(.A1(new_n580_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT118), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n843_), .B1(new_n854_), .B2(new_n857_), .ZN(G1340gat));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n638_), .B(new_n852_), .C1(new_n842_), .C2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n540_), .B2(G120gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n842_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n846_), .A2(KEYINPUT119), .A3(new_n638_), .A4(new_n852_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G120gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n842_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n835_), .A2(new_n841_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n790_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n632_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n631_), .A2(G127gat), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT120), .Z(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n853_), .B2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT121), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n853_), .B2(new_n688_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n646_), .A2(G134gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n873_), .B2(new_n880_), .ZN(G1343gat));
  INV_X1    g680(.A(new_n432_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n738_), .A2(new_n882_), .A3(new_n788_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n872_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n639_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n638_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n884_), .A2(new_n632_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n885_), .B2(new_n645_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n682_), .A2(G162gat), .A3(new_n685_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n885_), .B2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n635_), .A2(new_n338_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n738_), .A2(new_n273_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n849_), .B2(new_n841_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n311_), .B1(new_n898_), .B2(new_n639_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n901_));
  OR3_X1    g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n901_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT123), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n899_), .A2(new_n905_), .A3(new_n901_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n900_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n902_), .A2(new_n904_), .A3(new_n906_), .A4(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n291_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n898_), .A2(new_n639_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1348gat));
  AOI21_X1  g710(.A(G176gat), .B1(new_n898_), .B2(new_n638_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n845_), .A2(new_n272_), .ZN(new_n913_));
  AND4_X1   g712(.A1(G176gat), .A2(new_n738_), .A3(new_n638_), .A4(new_n896_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  INV_X1    g714(.A(new_n898_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n916_), .A2(new_n300_), .A3(new_n632_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n913_), .A2(new_n631_), .A3(new_n738_), .A4(new_n896_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n279_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n916_), .B2(new_n688_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n898_), .A2(new_n295_), .A3(new_n645_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  XOR2_X1   g721(.A(new_n922_), .B(KEYINPUT125), .Z(G1351gat));
  OR2_X1    g722(.A1(new_n249_), .A2(KEYINPUT127), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n249_), .A2(KEYINPUT127), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n702_), .A2(new_n450_), .A3(new_n882_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n872_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT126), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n872_), .A2(new_n929_), .A3(new_n926_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n924_), .B(new_n925_), .C1(new_n931_), .C2(new_n640_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n930_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n933_), .A2(KEYINPUT127), .A3(new_n249_), .A4(new_n639_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(G1352gat));
  OAI21_X1  g734(.A(G204gat), .B1(new_n931_), .B2(new_n540_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n246_), .A3(new_n638_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1353gat));
  OR2_X1    g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n933_), .B2(new_n631_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n931_), .A2(new_n632_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n931_), .B2(new_n688_), .ZN(new_n944_));
  INV_X1    g743(.A(G218gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n933_), .A2(new_n945_), .A3(new_n645_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1355gat));
endmodule


