//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n851_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  OR4_X1    g009(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n211_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(new_n222_), .B2(KEYINPUT66), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n214_), .A3(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n210_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n210_), .A2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n230_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n226_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n225_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G43gat), .B(G50gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  AOI211_X1 g042(.A(KEYINPUT72), .B(new_n208_), .C1(new_n240_), .C2(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n234_), .A2(new_n237_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  INV_X1    g045(.A(new_n239_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .A4(new_n226_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n238_), .B2(new_n239_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n243_), .B(KEYINPUT15), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n244_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n207_), .A3(new_n205_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n205_), .A2(new_n207_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n244_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G190gat), .B(G218gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G134gat), .B(G162gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT36), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(KEYINPUT36), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n262_), .A3(new_n255_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G231gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G57gat), .B(G64gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n280_));
  XOR2_X1   g079(.A(G71gat), .B(G78gat), .Z(new_n281_));
  OR2_X1    g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n279_), .A2(KEYINPUT11), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n282_), .B(KEYINPUT68), .C1(new_n283_), .C2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n278_), .B(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n291_));
  XOR2_X1   g090(.A(G127gat), .B(G155gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(G183gat), .B(G211gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n290_), .A2(new_n291_), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT76), .ZN(new_n299_));
  INV_X1    g098(.A(new_n278_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n300_), .A2(new_n285_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n285_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n202_), .B1(new_n269_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n240_), .B(new_n285_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G230gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT12), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n240_), .B2(new_n285_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n240_), .A2(new_n285_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n314_), .A2(new_n309_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT5), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G176gat), .B(G204gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n311_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT69), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n311_), .A2(new_n317_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n321_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(KEYINPUT69), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT13), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT13), .B1(new_n326_), .B2(new_n328_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n306_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n267_), .A2(new_n334_), .A3(KEYINPUT77), .A4(new_n268_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n307_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT78), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n250_), .A2(new_n276_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n276_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n243_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G229gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n276_), .B(new_n243_), .Z(new_n347_));
  AOI22_X1  g146(.A1(new_n340_), .A2(new_n346_), .B1(new_n347_), .B2(new_n345_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G141gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G169gat), .B(G197gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n348_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G218gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G211gat), .ZN(new_n355_));
  INV_X1    g154(.A(G211gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G218gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT87), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G197gat), .A2(G204gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT21), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT21), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n362_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n359_), .A2(new_n361_), .A3(new_n365_), .A4(new_n368_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n367_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n355_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n360_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI22_X1  g176(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n377_), .A2(new_n378_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G155gat), .ZN(new_n384_));
  INV_X1    g183(.A(G162gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT83), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(G155gat), .B2(G162gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT1), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n386_), .A2(new_n391_), .A3(new_n388_), .A4(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G141gat), .B(G148gat), .Z(new_n395_));
  AOI22_X1  g194(.A1(new_n383_), .A2(new_n390_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n374_), .B1(KEYINPUT29), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(G233gat), .B1(KEYINPUT86), .B2(G228gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(KEYINPUT86), .B2(G228gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n369_), .A2(new_n373_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(KEYINPUT85), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n398_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT88), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n397_), .A2(KEYINPUT29), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G22gat), .B(G50gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT28), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n403_), .A2(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n406_), .A2(new_n412_), .A3(new_n405_), .A4(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT22), .B(G169gat), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n420_), .A2(new_n421_), .B1(G169gat), .B2(G176gat), .ZN(new_n422_));
  INV_X1    g221(.A(G183gat), .ZN(new_n423_));
  INV_X1    g222(.A(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n425_), .B(new_n428_), .C1(new_n429_), .C2(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n422_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n426_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n427_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT26), .B(G190gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT25), .B1(new_n436_), .B2(new_n423_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT25), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT24), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(G169gat), .B2(G176gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n441_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n434_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n431_), .A2(new_n446_), .A3(new_n369_), .A4(new_n373_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT81), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT23), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n427_), .A2(KEYINPUT81), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n432_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n424_), .A2(KEYINPUT26), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT26), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G190gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n438_), .A2(G183gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n423_), .A2(KEYINPUT25), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n451_), .A2(new_n457_), .A3(new_n428_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n427_), .A2(KEYINPUT81), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n448_), .A2(KEYINPUT23), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n432_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n426_), .A2(KEYINPUT23), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n425_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n458_), .A2(new_n445_), .B1(new_n463_), .B2(new_n422_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n447_), .B(KEYINPUT20), .C1(new_n464_), .C2(new_n374_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G226gat), .A2(G233gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT19), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G64gat), .B(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n374_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n431_), .A2(new_n446_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n401_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n467_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n474_), .A2(new_n476_), .A3(KEYINPUT20), .A4(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n468_), .A2(new_n473_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n473_), .B1(new_n468_), .B2(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(KEYINPUT27), .ZN(new_n482_));
  INV_X1    g281(.A(new_n479_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n465_), .A2(new_n467_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n463_), .A2(new_n422_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n445_), .A2(new_n451_), .A3(new_n428_), .A4(new_n457_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT20), .B1(new_n487_), .B2(new_n401_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n488_), .A2(KEYINPUT96), .B1(new_n475_), .B2(new_n401_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n490_), .A3(KEYINPUT20), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n484_), .B1(new_n492_), .B2(new_n467_), .ZN(new_n493_));
  OAI211_X1 g292(.A(KEYINPUT27), .B(new_n483_), .C1(new_n493_), .C2(new_n473_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n482_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n417_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G127gat), .B(G134gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G120gat), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n498_), .A2(new_n499_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n502_), .A2(new_n396_), .A3(KEYINPUT4), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n383_), .A2(new_n390_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n394_), .A2(new_n395_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT90), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n502_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n500_), .A2(new_n501_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n396_), .A2(KEYINPUT90), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n506_), .B1(new_n513_), .B2(KEYINPUT4), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n515_));
  AOI211_X1 g314(.A(KEYINPUT91), .B(new_n515_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n505_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n504_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G1gat), .B(G29gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT92), .B(G85gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT0), .B(G57gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(new_n518_), .A3(new_n524_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G71gat), .B(G99gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G43gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n475_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n502_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G227gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(G15gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT30), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT31), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n533_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n497_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT97), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n473_), .A2(KEYINPUT32), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n493_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n477_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n546_));
  OAI211_X1 g345(.A(KEYINPUT97), .B(new_n545_), .C1(new_n546_), .C2(new_n484_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n468_), .A2(new_n478_), .A3(new_n543_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n517_), .A2(KEYINPUT33), .A3(new_n518_), .A4(new_n524_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n503_), .B1(G225gat), .B2(G233gat), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n504_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT94), .B1(new_n555_), .B2(new_n524_), .ZN(new_n556_));
  OR3_X1    g355(.A1(new_n555_), .A2(KEYINPUT94), .A3(new_n524_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n554_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n552_), .A2(new_n481_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n527_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n527_), .A2(KEYINPUT93), .A3(new_n560_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n559_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n551_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n552_), .A2(new_n481_), .A3(new_n558_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n564_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT93), .B1(new_n527_), .B2(new_n560_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n568_), .B(new_n566_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n416_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n414_), .A2(new_n529_), .A3(new_n415_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(new_n495_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n539_), .B1(new_n573_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n541_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT95), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n571_), .A3(new_n551_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n575_), .B1(new_n582_), .B2(new_n416_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT98), .B1(new_n583_), .B2(new_n539_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n353_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n337_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n337_), .A2(KEYINPUT99), .A3(new_n585_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n271_), .A3(new_n528_), .A4(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n264_), .B(KEYINPUT101), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n352_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT100), .B(new_n352_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n600_), .A3(new_n334_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n529_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n590_), .A2(new_n591_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n602_), .A3(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(new_n495_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(G8gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n588_), .A2(new_n589_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G8gat), .B1(new_n601_), .B2(new_n605_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT39), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n609_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(new_n539_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G15gat), .B1(new_n601_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT41), .Z(new_n618_));
  NAND4_X1  g417(.A1(new_n588_), .A2(new_n535_), .A3(new_n539_), .A4(new_n589_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1326gat));
  OAI21_X1  g419(.A(G22gat), .B1(new_n601_), .B2(new_n416_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT42), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n416_), .A2(G22gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n588_), .A2(new_n589_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(G1327gat));
  NOR2_X1   g424(.A1(new_n334_), .A2(new_n264_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n333_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n585_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(G29gat), .B1(new_n628_), .B2(new_n528_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  INV_X1    g429(.A(new_n269_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n579_), .B2(new_n584_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n630_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n580_), .A2(KEYINPUT95), .B1(new_n548_), .B2(new_n550_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n417_), .B1(new_n635_), .B2(new_n571_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n578_), .B(new_n616_), .C1(new_n636_), .C2(new_n575_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n541_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n577_), .A2(new_n578_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n269_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n634_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n598_), .A2(new_n306_), .A3(new_n599_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT104), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT44), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n648_), .B(new_n645_), .C1(new_n634_), .C2(new_n642_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n528_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n629_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  XNOR2_X1  g451(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G36gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n650_), .B2(new_n495_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n495_), .B(KEYINPUT106), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n628_), .A2(new_n655_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT45), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n654_), .B1(new_n656_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n643_), .A2(new_n646_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n648_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n643_), .A2(KEYINPUT44), .A3(new_n646_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n495_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n660_), .A3(new_n653_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n668_), .ZN(G1329gat));
  INV_X1    g468(.A(G43gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n628_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n616_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n664_), .A2(new_n665_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n539_), .A2(G43gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT47), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT47), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n677_), .B(new_n672_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1330gat));
  OR3_X1    g478(.A1(new_n671_), .A2(G50gat), .A3(new_n416_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n650_), .A2(new_n681_), .A3(new_n417_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n650_), .B2(new_n417_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1331gat));
  AOI211_X1 g484(.A(new_n352_), .B(new_n333_), .C1(new_n579_), .C2(new_n584_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n686_), .A2(new_n307_), .A3(new_n335_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n528_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT109), .ZN(new_n689_));
  INV_X1    g488(.A(new_n333_), .ZN(new_n690_));
  AND4_X1   g489(.A1(new_n353_), .A2(new_n595_), .A3(new_n690_), .A4(new_n334_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(G57gat), .A3(new_n528_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n691_), .B2(new_n658_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT48), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n687_), .A2(new_n694_), .A3(new_n658_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1333gat));
  INV_X1    g497(.A(G71gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n691_), .B2(new_n539_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT49), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n539_), .A2(new_n699_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT110), .Z(new_n703_));
  NAND2_X1  g502(.A1(new_n687_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1334gat));
  INV_X1    g504(.A(G78gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n691_), .B2(new_n417_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT50), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n687_), .A2(new_n706_), .A3(new_n417_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1335gat));
  NAND2_X1  g509(.A1(new_n686_), .A2(new_n626_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(new_n218_), .A3(new_n528_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n333_), .A2(new_n352_), .A3(new_n334_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT43), .B1(new_n641_), .B2(KEYINPUT105), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n584_), .A2(new_n638_), .A3(new_n637_), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n633_), .B(new_n630_), .C1(new_n716_), .C2(new_n269_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n643_), .A2(KEYINPUT111), .A3(new_n714_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n529_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n713_), .B1(new_n722_), .B2(new_n218_), .ZN(G1336gat));
  NAND3_X1  g522(.A1(new_n712_), .A2(new_n219_), .A3(new_n495_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n657_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(new_n219_), .ZN(G1337gat));
  AND4_X1   g525(.A1(new_n539_), .A2(new_n712_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n616_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n213_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n728_), .C1(new_n729_), .C2(new_n213_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n712_), .A2(new_n214_), .A3(new_n417_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n643_), .A2(new_n417_), .A3(new_n714_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G106gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT53), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT53), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n735_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1339gat));
  NOR3_X1   g543(.A1(new_n497_), .A2(new_n616_), .A3(new_n529_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT57), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n324_), .B(new_n327_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n347_), .A2(new_n344_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n351_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT117), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n343_), .A2(new_n344_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n340_), .A2(new_n753_), .B1(new_n751_), .B2(KEYINPUT117), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n752_), .A2(new_n754_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n748_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n314_), .A2(new_n316_), .A3(new_n315_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n310_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(new_n310_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n317_), .A2(new_n763_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n760_), .A2(new_n761_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n317_), .A2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n317_), .A2(new_n763_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(KEYINPUT113), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT115), .B(new_n321_), .C1(new_n765_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT116), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n352_), .A2(new_n323_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n321_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT115), .B1(new_n773_), .B2(KEYINPUT116), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n757_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n264_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT118), .B(new_n747_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n755_), .A2(new_n323_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n776_), .B2(KEYINPUT56), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n317_), .A2(new_n766_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n768_), .A2(KEYINPUT113), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n786_), .B(new_n787_), .C1(new_n761_), .C2(new_n760_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n773_), .B1(new_n788_), .B2(new_n321_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n773_), .A3(new_n321_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n776_), .A2(KEYINPUT56), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT58), .A4(new_n783_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n269_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n776_), .A2(new_n777_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n352_), .A3(new_n323_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n770_), .B2(new_n771_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n756_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT57), .A3(new_n264_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n781_), .A2(new_n794_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT57), .B1(new_n798_), .B2(new_n264_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(KEYINPUT118), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n306_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n333_), .A2(new_n353_), .A3(new_n631_), .A4(new_n334_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT54), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT54), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n746_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n790_), .A2(new_n269_), .A3(new_n793_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n801_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n747_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(KEYINPUT119), .A3(new_n794_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n815_), .A3(new_n799_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n807_), .B1(new_n816_), .B2(new_n306_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n745_), .A2(new_n810_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n809_), .A2(new_n810_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819_), .B2(new_n353_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n809_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n353_), .A2(G113gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  OAI21_X1  g622(.A(G120gat), .B1(new_n819_), .B2(new_n333_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n825_));
  AOI21_X1  g624(.A(G120gat), .B1(new_n690_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n825_), .B2(G120gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n809_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(KEYINPUT120), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1341gat));
  OAI21_X1  g632(.A(G127gat), .B1(new_n819_), .B2(new_n306_), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n821_), .A2(G127gat), .A3(new_n306_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1342gat));
  OAI21_X1  g639(.A(G134gat), .B1(new_n819_), .B2(new_n631_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n593_), .A2(G134gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n821_), .B2(new_n842_), .ZN(G1343gat));
  AND2_X1   g642(.A1(new_n803_), .A2(new_n808_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n539_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n658_), .A2(new_n529_), .A3(new_n416_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n352_), .A3(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n846_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n333_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT122), .B(G148gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1345gat));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n306_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT61), .B(G155gat), .Z(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1346gat));
  OAI21_X1  g654(.A(G162gat), .B1(new_n849_), .B2(new_n631_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n594_), .A2(new_n385_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n849_), .B2(new_n857_), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n817_), .A2(new_n417_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n657_), .A2(new_n540_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n352_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G169gat), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n421_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n864_), .B(new_n865_), .C1(new_n866_), .C2(new_n861_), .ZN(G1348gat));
  NAND3_X1  g666(.A1(new_n859_), .A2(new_n690_), .A3(new_n860_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n844_), .A2(new_n417_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n690_), .A2(G176gat), .A3(new_n860_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n868_), .A2(new_n420_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  NAND2_X1  g670(.A1(new_n860_), .A2(new_n334_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n859_), .A2(new_n873_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n844_), .A2(new_n417_), .A3(new_n872_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G183gat), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1350gat));
  NAND4_X1  g677(.A1(new_n859_), .A2(new_n435_), .A3(new_n594_), .A4(new_n860_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n859_), .A2(new_n269_), .A3(new_n860_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n880_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT124), .B1(new_n880_), .B2(G190gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n879_), .B1(new_n881_), .B2(new_n882_), .ZN(G1351gat));
  NOR2_X1   g682(.A1(new_n657_), .A2(new_n574_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n845_), .A2(new_n352_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  OR2_X1    g685(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n845_), .A2(new_n884_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n333_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT126), .Z(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n887_), .B(new_n891_), .C1(new_n888_), .C2(new_n333_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1353gat));
  AND2_X1   g694(.A1(new_n845_), .A2(new_n884_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT63), .B(G211gat), .Z(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n334_), .A3(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n888_), .B2(new_n306_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1354gat));
  AOI21_X1  g700(.A(G218gat), .B1(new_n896_), .B2(new_n594_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n269_), .A2(G218gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT127), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n896_), .B2(new_n904_), .ZN(G1355gat));
endmodule


