//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT81), .B(G113gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G120gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n202_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT31), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n205_), .A2(new_n209_), .A3(KEYINPUT31), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT80), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT30), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AOI211_X1 g015(.A(KEYINPUT80), .B(KEYINPUT30), .C1(new_n212_), .C2(new_n213_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT77), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT78), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT78), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n222_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n221_), .B1(new_n232_), .B2(KEYINPUT24), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(KEYINPUT76), .A2(G190gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT26), .Z(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G183gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT75), .B(G183gat), .Z(new_n240_));
  OAI211_X1 g039(.A(new_n237_), .B(new_n239_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n233_), .A2(new_n235_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n220_), .B1(G190gat), .B2(new_n240_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G169gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n222_), .B1(new_n244_), .B2(new_n224_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(G71gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n218_), .A2(new_n253_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n251_), .B(new_n252_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G15gat), .B(G43gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT79), .B(G99gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(new_n259_), .A3(new_n255_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NOR4_X1   g065(.A1(KEYINPUT84), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT2), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n266_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n265_), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n276_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT83), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n279_), .A2(new_n284_), .A3(new_n276_), .A4(new_n280_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n273_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(new_n269_), .ZN(new_n288_));
  AOI221_X4 g087(.A(new_n264_), .B1(new_n275_), .B2(new_n276_), .C1(new_n286_), .C2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n288_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n275_), .A2(new_n276_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT85), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT29), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT88), .B(G197gat), .ZN(new_n295_));
  OAI211_X1 g094(.A(KEYINPUT21), .B(new_n294_), .C1(new_n295_), .C2(G204gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G197gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n296_), .B(new_n297_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n297_), .A2(KEYINPUT90), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(KEYINPUT90), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(new_n300_), .A3(KEYINPUT21), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT87), .B(G233gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT86), .B(G228gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n293_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n306_), .B(KEYINPUT91), .Z(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G78gat), .B(G106gat), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n311_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n289_), .A2(new_n292_), .A3(KEYINPUT29), .ZN(new_n321_));
  XOR2_X1   g120(.A(G22gat), .B(G50gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT28), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n319_), .A2(KEYINPUT92), .A3(new_n320_), .A4(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n320_), .A2(new_n327_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n328_), .A2(new_n324_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n263_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n210_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT96), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n290_), .A2(new_n205_), .A3(new_n209_), .A4(new_n291_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT96), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n335_), .B(new_n210_), .C1(new_n289_), .C2(new_n292_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .A4(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n331_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(KEYINPUT4), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n337_), .B1(new_n341_), .B2(new_n333_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G85gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT0), .B(G57gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n346_), .B(new_n337_), .C1(new_n341_), .C2(new_n333_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n330_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n328_), .A2(new_n324_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n319_), .A2(new_n320_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n353_), .A2(new_n325_), .A3(new_n262_), .A4(new_n261_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n306_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n242_), .A2(new_n355_), .A3(new_n246_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(new_n245_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n228_), .A2(new_n234_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n238_), .A2(G183gat), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(new_n239_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n233_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT93), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n233_), .A2(new_n366_), .A3(new_n359_), .A4(new_n363_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n358_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n356_), .B(KEYINPUT20), .C1(new_n368_), .C2(new_n355_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n355_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n371_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n247_), .B2(new_n306_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G8gat), .B(G36gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT95), .ZN(new_n379_));
  XOR2_X1   g178(.A(G64gat), .B(G92gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n372_), .A2(new_n377_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT99), .ZN(new_n386_));
  INV_X1    g185(.A(new_n358_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n312_), .A2(new_n364_), .A3(new_n387_), .ZN(new_n388_));
  AOI211_X1 g187(.A(new_n386_), .B(new_n374_), .C1(new_n388_), .C2(new_n376_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT99), .B1(new_n369_), .B2(new_n371_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n376_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n371_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n389_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT27), .B(new_n385_), .C1(new_n393_), .C2(new_n384_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT27), .ZN(new_n395_));
  INV_X1    g194(.A(new_n385_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n384_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n354_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n350_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n349_), .A2(KEYINPUT97), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT33), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n396_), .A2(new_n397_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n340_), .A2(KEYINPUT4), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT98), .B(new_n333_), .C1(new_n404_), .C2(new_n339_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n340_), .A2(new_n333_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(new_n346_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT98), .ZN(new_n408_));
  INV_X1    g207(.A(new_n333_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n341_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n349_), .A2(KEYINPUT97), .A3(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n402_), .A2(new_n403_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n372_), .A2(new_n377_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n384_), .A2(KEYINPUT32), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n416_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n393_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n414_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n354_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n400_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G85gat), .B(G92gat), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT9), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT10), .B(G99gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT64), .B(G106gat), .ZN(new_n429_));
  OAI221_X1 g228(.A(new_n426_), .B1(KEYINPUT9), .B2(new_n427_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  OR3_X1    g229(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n430_), .B1(KEYINPUT8), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT6), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n425_), .A2(KEYINPUT8), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n433_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n436_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT8), .A3(new_n425_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G29gat), .B(G36gat), .ZN(new_n444_));
  INV_X1    g243(.A(G50gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT68), .B(G43gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n448_), .B(KEYINPUT15), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n443_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G232gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT35), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT69), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n451_), .A2(KEYINPUT69), .A3(new_n443_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n450_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT35), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n455_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n457_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G190gat), .B(G218gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G134gat), .B(G162gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(KEYINPUT70), .B2(KEYINPUT36), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n464_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n467_), .B(KEYINPUT36), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n464_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n475_), .A3(KEYINPUT37), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT71), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n464_), .A2(KEYINPUT71), .A3(new_n474_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n472_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n476_), .B1(new_n480_), .B2(KEYINPUT37), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G78gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT11), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(KEYINPUT11), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n482_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G231gat), .A2(G233gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491_));
  INV_X1    g290(.A(G1gat), .ZN(new_n492_));
  INV_X1    g291(.A(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G8gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT72), .Z(new_n498_));
  XNOR2_X1  g297(.A(new_n490_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT73), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G127gat), .B(G155gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(G211gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT16), .B(G183gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n501_), .B(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(new_n506_), .A3(new_n505_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n424_), .A2(new_n481_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n488_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n443_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n437_), .A2(new_n438_), .A3(new_n442_), .A4(new_n488_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(KEYINPUT12), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT12), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n443_), .A2(new_n517_), .A3(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n515_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT5), .B(G176gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G204gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n521_), .A2(new_n524_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT13), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n449_), .A2(new_n497_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n451_), .B2(new_n497_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT74), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n448_), .B(new_n497_), .Z(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(G229gat), .A3(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n512_), .A2(new_n536_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n348_), .A2(new_n349_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n492_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT38), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT100), .ZN(new_n557_));
  INV_X1    g356(.A(new_n534_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n551_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n424_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n480_), .A2(new_n511_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n492_), .B1(new_n563_), .B2(new_n553_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n555_), .B2(new_n554_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(new_n565_), .ZN(G1324gat));
  NAND2_X1  g365(.A1(new_n394_), .A2(new_n398_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G8gat), .B1(new_n562_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT39), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n552_), .A2(new_n493_), .A3(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT40), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(G1325gat));
  INV_X1    g373(.A(G15gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n563_), .B2(new_n263_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT41), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n552_), .A2(new_n575_), .A3(new_n263_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1326gat));
  NAND2_X1  g378(.A1(new_n353_), .A2(new_n325_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(G22gat), .B1(new_n562_), .B2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT101), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT42), .ZN(new_n584_));
  INV_X1    g383(.A(G22gat), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n552_), .A2(new_n585_), .A3(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(G1327gat));
  NAND2_X1  g386(.A1(new_n480_), .A2(new_n511_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n560_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(G29gat), .B1(new_n591_), .B2(new_n553_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT43), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT102), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n354_), .B1(new_n414_), .B2(new_n421_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n481_), .B(new_n594_), .C1(new_n595_), .C2(new_n400_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n511_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n350_), .A2(new_n399_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n349_), .A2(KEYINPUT97), .A3(new_n412_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n412_), .B1(new_n349_), .B2(KEYINPUT97), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n411_), .A2(new_n403_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n603_), .A2(new_n604_), .B1(new_n420_), .B2(new_n418_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n605_), .B2(new_n354_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n599_), .B1(new_n606_), .B2(new_n481_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n597_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n558_), .A2(new_n559_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n608_), .A2(KEYINPUT44), .A3(new_n609_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n612_), .A2(new_n553_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n592_), .B1(new_n614_), .B2(G29gat), .ZN(G1328gat));
  XOR2_X1   g414(.A(new_n567_), .B(KEYINPUT103), .Z(new_n616_));
  NOR3_X1   g415(.A1(new_n590_), .A2(G36gat), .A3(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT45), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n567_), .A3(new_n613_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G36gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n620_), .A3(KEYINPUT46), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1329gat));
  NAND4_X1  g424(.A1(new_n612_), .A2(G43gat), .A3(new_n263_), .A4(new_n613_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n590_), .B1(new_n262_), .B2(new_n261_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(G43gat), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g428(.A1(new_n612_), .A2(new_n580_), .A3(new_n613_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G50gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n591_), .A2(new_n445_), .A3(new_n580_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT104), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n631_), .A2(new_n635_), .A3(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(G1331gat));
  NOR2_X1   g436(.A1(new_n534_), .A2(new_n551_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n512_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n553_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(G57gat), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n536_), .A2(new_n424_), .A3(new_n551_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n561_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n553_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n642_), .B1(G57gat), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT105), .ZN(G1332gat));
  OAI21_X1  g447(.A(G64gat), .B1(new_n644_), .B2(new_n616_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT106), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT48), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n639_), .A2(G64gat), .A3(new_n616_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(G1333gat));
  AOI21_X1  g454(.A(new_n249_), .B1(new_n645_), .B2(new_n263_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n640_), .A2(new_n249_), .A3(new_n263_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1334gat));
  OR3_X1    g459(.A1(new_n639_), .A2(G78gat), .A3(new_n581_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n645_), .A2(new_n580_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(G78gat), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n662_), .B2(G78gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1335gat));
  NAND2_X1  g468(.A1(new_n643_), .A2(new_n589_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G85gat), .B1(new_n671_), .B2(new_n553_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n481_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n598_), .B1(new_n424_), .B2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n511_), .A3(new_n596_), .A4(new_n638_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n672_), .B1(new_n676_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g476(.A(G92gat), .B1(new_n671_), .B2(new_n567_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n675_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(G92gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n616_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1337gat));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n263_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G99gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n428_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n671_), .A2(new_n685_), .A3(new_n263_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n608_), .A2(new_n689_), .A3(new_n580_), .A4(new_n638_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT110), .B1(new_n675_), .B2(new_n581_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(G106gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT52), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT52), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n690_), .A2(new_n691_), .A3(new_n694_), .A4(G106gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n670_), .A2(new_n429_), .A3(new_n581_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT53), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n696_), .A2(new_n700_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1339gat));
  INV_X1    g501(.A(G113gat), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n568_), .A2(new_n553_), .A3(new_n263_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n542_), .A2(new_n540_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n538_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n547_), .B(new_n705_), .C1(new_n706_), .C2(new_n540_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n550_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n532_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT55), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n521_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n516_), .A2(new_n523_), .A3(new_n518_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n519_), .A2(KEYINPUT55), .A3(new_n520_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT56), .B1(new_n714_), .B2(new_n529_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n709_), .B1(new_n715_), .B2(KEYINPUT112), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n529_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n714_), .A2(KEYINPUT56), .A3(new_n529_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n708_), .B(new_n716_), .C1(new_n721_), .C2(KEYINPUT112), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT58), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT58), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(new_n723_), .A3(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n481_), .A3(new_n727_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n551_), .A2(KEYINPUT111), .A3(new_n532_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT111), .B1(new_n551_), .B2(new_n532_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n721_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n533_), .A2(new_n708_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n480_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT57), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n737_), .B(new_n480_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n510_), .B1(new_n728_), .B2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n673_), .A2(new_n534_), .A3(new_n510_), .A4(new_n559_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n581_), .B(new_n704_), .C1(new_n740_), .C2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n703_), .B1(new_n744_), .B2(new_n559_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n744_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT59), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n744_), .A2(KEYINPUT59), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT115), .B(G113gat), .Z(new_n752_));
  NAND4_X1  g551(.A1(new_n750_), .A2(new_n551_), .A3(new_n751_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n745_), .A2(new_n746_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n747_), .A2(new_n753_), .A3(new_n754_), .ZN(G1340gat));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n751_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G120gat), .B1(new_n756_), .B2(new_n536_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n206_), .B1(new_n534_), .B2(KEYINPUT60), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n748_), .B(new_n758_), .C1(KEYINPUT60), .C2(new_n206_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1341gat));
  AOI21_X1  g559(.A(G127gat), .B1(new_n748_), .B2(new_n510_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n756_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n510_), .A2(G127gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(G1342gat));
  AOI21_X1  g563(.A(G134gat), .B1(new_n748_), .B2(new_n480_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT116), .B(G134gat), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n673_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n762_), .B2(new_n767_), .ZN(G1343gat));
  NOR2_X1   g567(.A1(new_n581_), .A2(new_n263_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n553_), .B(new_n769_), .C1(new_n740_), .C2(new_n743_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(new_n681_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n551_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g572(.A(new_n536_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT117), .B(G148gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(G1345gat));
  XNOR2_X1  g576(.A(KEYINPUT61), .B(G155gat), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  XOR2_X1   g578(.A(KEYINPUT118), .B(KEYINPUT119), .Z(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n771_), .B2(new_n510_), .ZN(new_n782_));
  NOR4_X1   g581(.A1(new_n770_), .A2(new_n511_), .A3(new_n681_), .A4(new_n780_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n769_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n722_), .A2(new_n723_), .A3(new_n726_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n726_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n673_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n734_), .A2(new_n735_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n737_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n734_), .A2(KEYINPUT57), .A3(new_n735_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n511_), .B1(new_n788_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n741_), .B(KEYINPUT54), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n785_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n553_), .A3(new_n616_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n780_), .B1(new_n796_), .B2(new_n511_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n771_), .A2(new_n510_), .A3(new_n781_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n778_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n784_), .A2(new_n799_), .ZN(G1346gat));
  INV_X1    g599(.A(G162gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n771_), .B2(new_n481_), .ZN(new_n802_));
  NOR4_X1   g601(.A1(new_n770_), .A2(G162gat), .A3(new_n735_), .A4(new_n681_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT120), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G162gat), .B1(new_n796_), .B2(new_n673_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n771_), .A2(new_n801_), .A3(new_n480_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(G1347gat));
  NOR2_X1   g608(.A1(new_n616_), .A2(new_n553_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(new_n263_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n581_), .B(new_n811_), .C1(new_n740_), .C2(new_n743_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT121), .B1(new_n812_), .B2(new_n559_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n580_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n551_), .A4(new_n811_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n813_), .A2(new_n816_), .A3(G169gat), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n812_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n244_), .A3(new_n551_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n813_), .A2(new_n816_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(G1348gat));
  AOI21_X1  g622(.A(G176gat), .B1(new_n820_), .B2(new_n558_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n814_), .A2(KEYINPUT122), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n581_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AND4_X1   g627(.A1(new_n774_), .A2(new_n825_), .A3(new_n811_), .A4(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n829_), .B2(G176gat), .ZN(G1349gat));
  INV_X1    g629(.A(new_n361_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n814_), .A2(new_n510_), .A3(new_n831_), .A4(new_n811_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT123), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n820_), .A2(new_n834_), .A3(new_n510_), .A4(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n240_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n825_), .A2(new_n828_), .A3(new_n510_), .A4(new_n811_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1350gat));
  OAI21_X1  g638(.A(G190gat), .B1(new_n812_), .B2(new_n673_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n480_), .A2(new_n362_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n812_), .B2(new_n841_), .ZN(G1351gat));
  NAND2_X1  g641(.A1(new_n795_), .A2(new_n810_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n551_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n536_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(new_n298_), .ZN(G1353gat));
  AOI21_X1  g647(.A(new_n511_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT124), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(KEYINPUT124), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n843_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1354gat));
  XOR2_X1   g654(.A(KEYINPUT125), .B(G218gat), .Z(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n844_), .B2(new_n480_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n481_), .A2(new_n856_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT126), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n844_), .B2(new_n859_), .ZN(G1355gat));
endmodule


