//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  NAND2_X1  g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(G106gat), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(KEYINPUT9), .B2(new_n202_), .ZN(new_n215_));
  OR3_X1    g014(.A1(new_n208_), .A2(new_n209_), .A3(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n209_), .B1(new_n208_), .B2(new_n215_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G57gat), .B(G64gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(KEYINPUT11), .ZN(new_n222_));
  XOR2_X1   g021(.A(G71gat), .B(G78gat), .Z(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n222_), .A2(new_n223_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n214_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT7), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT65), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n227_), .B1(new_n233_), .B2(new_n205_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT66), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n214_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT8), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(new_n234_), .B2(KEYINPUT66), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n219_), .B(new_n226_), .C1(new_n236_), .C2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n218_), .B1(new_n242_), .B2(new_n235_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(KEYINPUT67), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n224_), .A2(new_n245_), .A3(new_n225_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n219_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n226_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT12), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G230gat), .A2(G233gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n243_), .A2(new_n226_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n241_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT69), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n254_), .A2(new_n258_), .A3(new_n265_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(KEYINPUT13), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT71), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT71), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G1gat), .B(G8gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT72), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT72), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(G231gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n244_), .A2(new_n246_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G127gat), .B(G155gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT16), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT17), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n294_), .A2(new_n295_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n226_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n291_), .A2(new_n250_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n299_), .B(KEYINPUT17), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT73), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G29gat), .B(G36gat), .Z(new_n310_));
  XOR2_X1   g109(.A(G43gat), .B(G50gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT15), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n249_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n243_), .A2(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT34), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n317_), .A2(KEYINPUT35), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n314_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(KEYINPUT35), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G190gat), .B(G218gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G134gat), .B(G162gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT36), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(KEYINPUT35), .A3(new_n317_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n321_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n324_), .B(KEYINPUT36), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n321_), .B2(new_n326_), .ZN(new_n330_));
  OR3_X1    g129(.A1(new_n327_), .A2(new_n330_), .A3(KEYINPUT37), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT37), .B1(new_n327_), .B2(new_n330_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n277_), .A2(new_n309_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(KEYINPUT24), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n347_), .B1(new_n350_), .B2(KEYINPUT24), .ZN(new_n351_));
  OR2_X1    g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n341_), .A2(new_n352_), .A3(new_n342_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n353_), .A2(new_n348_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT22), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(G169gat), .ZN(new_n356_));
  INV_X1    g155(.A(G169gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(KEYINPUT22), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT75), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT76), .B(G176gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(KEYINPUT22), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n344_), .A2(new_n351_), .B1(new_n354_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366_));
  INV_X1    g165(.A(G43gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n365_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G15gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT30), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n373_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G127gat), .B(G134gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT77), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT31), .ZN(new_n381_));
  AND4_X1   g180(.A1(KEYINPUT78), .A2(new_n374_), .A3(new_n375_), .A4(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT78), .B1(new_n374_), .B2(new_n375_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n381_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(KEYINPUT78), .A3(new_n375_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n382_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G141gat), .A2(G148gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT79), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G141gat), .ZN(new_n393_));
  INV_X1    g192(.A(G148gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT1), .ZN(new_n398_));
  INV_X1    g197(.A(G155gat), .ZN(new_n399_));
  INV_X1    g198(.A(G162gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT80), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n401_), .A2(new_n403_), .B1(KEYINPUT1), .B2(new_n397_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n398_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n397_), .A2(KEYINPUT1), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT81), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n396_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n397_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415_));
  OAI22_X1  g214(.A1(new_n413_), .A2(new_n414_), .B1(new_n388_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(KEYINPUT2), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n392_), .B2(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT82), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n412_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n411_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  XOR2_X1   g222(.A(G22gat), .B(G50gat), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(new_n423_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n424_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n428_), .B1(new_n433_), .B2(new_n426_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n387_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n429_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n428_), .A3(new_n426_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(KEYINPUT91), .A3(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G78gat), .B(G106gat), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n441_), .B(KEYINPUT85), .Z(new_n442_));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n443_));
  INV_X1    g242(.A(G211gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(G218gat), .ZN(new_n445_));
  INV_X1    g244(.A(G218gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(G211gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n443_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G197gat), .A2(G204gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G197gat), .A2(G204gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT21), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(G211gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n444_), .A2(G218gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT87), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT87), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT87), .B1(new_n454_), .B2(new_n455_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n451_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT21), .A3(new_n449_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n452_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n457_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT88), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n462_), .B(new_n463_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n468_), .B2(new_n457_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n464_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n448_), .A2(new_n456_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT88), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT90), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n396_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n407_), .A2(new_n405_), .A3(new_n408_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n398_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n404_), .A2(new_n405_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n412_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n416_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n388_), .B(new_n389_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n417_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n419_), .B(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n483_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n423_), .B1(new_n482_), .B2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n471_), .B(new_n476_), .C1(new_n491_), .C2(KEYINPUT89), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT89), .B(KEYINPUT29), .C1(new_n411_), .C2(new_n421_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n442_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n442_), .B(KEYINPUT86), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(new_n491_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n440_), .B1(new_n495_), .B2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT29), .B1(new_n411_), .B2(new_n421_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n503_), .A2(new_n493_), .A3(new_n476_), .A4(new_n471_), .ZN(new_n504_));
  AOI211_X1 g303(.A(new_n498_), .B(new_n439_), .C1(new_n504_), .C2(new_n442_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n435_), .B(new_n438_), .C1(new_n500_), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n495_), .A2(new_n499_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n439_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT91), .B1(new_n436_), .B2(new_n437_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n495_), .A2(new_n499_), .A3(new_n440_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G1gat), .B(G29gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G85gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n377_), .B(new_n378_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n411_), .B2(new_n421_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n422_), .A2(new_n380_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G225gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n517_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT99), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT99), .B(new_n517_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT4), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n422_), .A2(new_n380_), .A3(KEYINPUT4), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n523_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n532_), .A3(new_n524_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n517_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n519_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT93), .B1(new_n356_), .B2(new_n358_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n355_), .A2(G169gat), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n361_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n360_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n353_), .A2(KEYINPUT94), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n341_), .A2(new_n352_), .A3(new_n548_), .A4(new_n342_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n546_), .A2(new_n547_), .A3(new_n348_), .A4(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n349_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n345_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n338_), .A3(new_n343_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n466_), .A2(new_n365_), .A3(new_n470_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT20), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G226gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT19), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G8gat), .B(G36gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT18), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G64gat), .B(G92gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n466_), .A2(new_n470_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n555_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n555_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n472_), .A2(new_n475_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(KEYINPUT95), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n560_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT20), .B(new_n573_), .C1(new_n570_), .C2(new_n365_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n561_), .B(new_n565_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT96), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n577_));
  INV_X1    g376(.A(new_n365_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n567_), .B2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n568_), .A2(new_n579_), .A3(new_n573_), .A4(new_n571_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n561_), .A4(new_n565_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n561_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n565_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n541_), .A2(new_n576_), .A3(new_n582_), .A4(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n539_), .A2(new_n540_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n535_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n565_), .A2(KEYINPUT32), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n561_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n471_), .A2(new_n476_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n569_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n573_), .B1(new_n592_), .B2(new_n579_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n558_), .A2(new_n560_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n590_), .B1(new_n595_), .B2(new_n589_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n537_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n539_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n539_), .A2(KEYINPUT100), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n596_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n512_), .B1(new_n588_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n512_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n599_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n597_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n605_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n576_), .A2(new_n585_), .A3(new_n582_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT27), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n584_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n575_), .A2(KEYINPUT27), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n608_), .A2(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n386_), .B1(new_n603_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(new_n386_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n612_), .A2(KEYINPUT101), .A3(new_n512_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT101), .B1(new_n612_), .B2(new_n512_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n608_), .A2(new_n609_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n611_), .A2(new_n610_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n512_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n612_), .A2(KEYINPUT101), .A3(new_n512_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT102), .A3(new_n616_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n614_), .B1(new_n621_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n289_), .B(new_n312_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(G229gat), .A3(G233gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n313_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n289_), .A2(new_n312_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT74), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n638_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n637_), .A3(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n630_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n335_), .A2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT103), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n605_), .A2(new_n601_), .A3(new_n606_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n283_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n277_), .A2(new_n646_), .A3(new_n309_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n327_), .A2(new_n330_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n630_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n607_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n651_), .A2(new_n652_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n658_), .A3(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(new_n612_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n649_), .A2(new_n284_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n657_), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT39), .B(new_n284_), .C1(new_n663_), .C2(new_n661_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n661_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G8gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n662_), .B(KEYINPUT40), .C1(new_n667_), .C2(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(new_n386_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G15gat), .B1(new_n657_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT41), .Z(new_n675_));
  INV_X1    g474(.A(new_n648_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n371_), .A3(new_n386_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n657_), .B2(new_n512_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT42), .Z(new_n680_));
  NOR3_X1   g479(.A1(new_n648_), .A2(G22gat), .A3(new_n512_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  AND2_X1   g481(.A1(new_n275_), .A2(new_n276_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n647_), .A2(new_n683_), .A3(new_n309_), .A4(new_n655_), .ZN(new_n684_));
  INV_X1    g483(.A(G29gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n650_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n333_), .B2(KEYINPUT104), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n630_), .B2(new_n333_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n586_), .A2(new_n587_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n534_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n602_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n604_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n613_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n673_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT102), .B1(new_n628_), .B2(new_n616_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n620_), .B(new_n615_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n334_), .A3(new_n688_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n690_), .A2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n277_), .A2(new_n646_), .A3(new_n308_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n701_), .B2(new_n702_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n650_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n687_), .B1(new_n707_), .B2(G29gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT105), .B(new_n685_), .C1(new_n706_), .C2(new_n650_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n686_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  NOR3_X1   g509(.A1(new_n704_), .A2(new_n705_), .A3(new_n612_), .ZN(new_n711_));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n684_), .A2(new_n712_), .A3(new_n661_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  OR3_X1    g516(.A1(new_n713_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n713_), .B2(new_n716_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1329gat));
  NAND3_X1  g519(.A1(new_n706_), .A2(G43gat), .A3(new_n386_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n684_), .A2(new_n386_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n367_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n684_), .A2(new_n727_), .A3(new_n604_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n630_), .A2(new_n689_), .A3(new_n333_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n688_), .B1(new_n699_), .B2(new_n334_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n702_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n604_), .A3(new_n703_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G50gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n728_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT109), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(new_n728_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1331gat));
  AND4_X1   g541(.A1(new_n646_), .A2(new_n656_), .A3(new_n277_), .A4(new_n308_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(G57gat), .A3(new_n650_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT110), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(KEYINPUT110), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n334_), .A2(new_n309_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n277_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n630_), .A2(new_n645_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n650_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n745_), .A2(new_n746_), .A3(new_n752_), .ZN(G1332gat));
  INV_X1    g552(.A(G64gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n754_), .A3(new_n661_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n743_), .A2(new_n661_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(G64gat), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT48), .B(new_n754_), .C1(new_n743_), .C2(new_n661_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT111), .ZN(G1333gat));
  NAND2_X1  g560(.A1(new_n743_), .A2(new_n386_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G71gat), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT49), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n673_), .A2(G71gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT112), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n750_), .B2(new_n766_), .ZN(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n743_), .B2(new_n604_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n751_), .A2(new_n768_), .A3(new_n604_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n701_), .B(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n683_), .A2(new_n645_), .A3(new_n308_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776_), .B2(new_n607_), .ZN(new_n777_));
  AND4_X1   g576(.A1(new_n277_), .A2(new_n749_), .A3(new_n309_), .A4(new_n655_), .ZN(new_n778_));
  INV_X1    g577(.A(G85gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n650_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n776_), .B2(new_n612_), .ZN(new_n782_));
  INV_X1    g581(.A(G92gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n778_), .A2(new_n783_), .A3(new_n661_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n776_), .B2(new_n673_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n673_), .A2(new_n207_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n778_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT51), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(new_n791_), .A3(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1338gat));
  INV_X1    g592(.A(G106gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n778_), .A2(new_n794_), .A3(new_n604_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n775_), .A2(new_n701_), .A3(new_n604_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(G106gat), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT52), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(KEYINPUT52), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n631_), .A2(new_n636_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n636_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n633_), .A2(new_n634_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n642_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n644_), .A2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT118), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n269_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n242_), .A2(new_n235_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n247_), .B1(new_n810_), .B2(new_n219_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n257_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT12), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n243_), .B2(new_n226_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n812_), .A2(KEYINPUT55), .A3(new_n253_), .A4(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n814_), .B(new_n241_), .C1(new_n243_), .C2(new_n247_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n255_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n252_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n253_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n255_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n817_), .A2(new_n820_), .A3(new_n821_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n266_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT116), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n823_), .A2(KEYINPUT116), .A3(new_n825_), .A4(new_n266_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n268_), .A2(new_n645_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n809_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n827_), .A2(KEYINPUT117), .A3(new_n828_), .A4(new_n829_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n655_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n268_), .B(new_n808_), .C1(new_n824_), .C2(KEYINPUT56), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n825_), .B1(new_n823_), .B2(new_n266_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n334_), .ZN(new_n840_));
  OAI22_X1  g639(.A1(new_n834_), .A2(KEYINPUT57), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n842_), .B(new_n655_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n309_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n747_), .A2(new_n646_), .A3(new_n274_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT54), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n628_), .A2(new_n650_), .A3(new_n386_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT119), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n802_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n849_), .B(new_n853_), .C1(new_n844_), .C2(new_n846_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT121), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n850_), .A3(new_n852_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n849_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n856_), .B(new_n857_), .C1(new_n802_), .C2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n645_), .A2(KEYINPUT122), .A3(G113gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(KEYINPUT122), .B2(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G113gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n858_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n646_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1340gat));
  XOR2_X1   g665(.A(KEYINPUT123), .B(G120gat), .Z(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n858_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n867_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n851_), .A2(new_n854_), .A3(new_n683_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n309_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n855_), .A2(new_n859_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n864_), .B2(new_n309_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1342gat));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n333_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n855_), .A2(new_n859_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n655_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n877_), .B1(new_n864_), .B2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1343gat));
  NOR4_X1   g681(.A1(new_n661_), .A2(new_n607_), .A3(new_n512_), .A4(new_n386_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n847_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n646_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n393_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n683_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n394_), .ZN(G1345gat));
  OAI21_X1  g687(.A(KEYINPUT124), .B1(new_n884_), .B2(new_n309_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n847_), .A2(new_n890_), .A3(new_n308_), .A4(new_n883_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n889_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n884_), .B2(new_n333_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n655_), .A2(new_n400_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n884_), .B2(new_n897_), .ZN(G1347gat));
  NAND3_X1  g697(.A1(new_n616_), .A2(new_n512_), .A3(new_n661_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n900_), .A2(new_n645_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n357_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n901_), .B2(new_n357_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n901_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(G1348gat));
  AND3_X1   g705(.A1(new_n900_), .A2(G176gat), .A3(new_n277_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n900_), .A2(new_n277_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n360_), .B2(new_n908_), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n900_), .A2(new_n308_), .ZN(new_n910_));
  MUX2_X1   g709(.A(new_n336_), .B(G183gat), .S(new_n910_), .Z(G1350gat));
  NAND3_X1  g710(.A1(new_n900_), .A2(new_n337_), .A3(new_n655_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n900_), .A2(new_n334_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n913_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT125), .B1(new_n913_), .B2(G190gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n912_), .B1(new_n914_), .B2(new_n915_), .ZN(G1351gat));
  NOR4_X1   g715(.A1(new_n612_), .A2(new_n512_), .A3(new_n650_), .A4(new_n386_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n847_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT126), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n847_), .A2(new_n920_), .A3(new_n917_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G197gat), .B1(new_n922_), .B2(new_n645_), .ZN(new_n923_));
  INV_X1    g722(.A(G197gat), .ZN(new_n924_));
  AOI211_X1 g723(.A(new_n924_), .B(new_n646_), .C1(new_n919_), .C2(new_n921_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1352gat));
  INV_X1    g725(.A(new_n921_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n920_), .B1(new_n847_), .B2(new_n917_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n277_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G204gat), .ZN(new_n930_));
  INV_X1    g729(.A(G204gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n922_), .A2(new_n931_), .A3(new_n277_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1353gat));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n309_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n922_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  AOI211_X1 g737(.A(new_n934_), .B(new_n938_), .C1(new_n919_), .C2(new_n921_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1354gat));
  NAND2_X1  g739(.A1(new_n922_), .A2(new_n655_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT127), .B(G218gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n333_), .A2(new_n942_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n941_), .A2(new_n942_), .B1(new_n922_), .B2(new_n943_), .ZN(G1355gat));
endmodule


