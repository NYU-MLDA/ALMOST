//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G197gat), .B2(G204gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n202_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(G197gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n203_), .A2(new_n205_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n210_), .C1(new_n211_), .C2(new_n204_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n210_), .B1(new_n211_), .B2(new_n204_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(new_n207_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n219_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT93), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI211_X1 g025(.A(KEYINPUT93), .B(new_n219_), .C1(new_n221_), .C2(new_n223_), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  INV_X1    g030(.A(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n226_), .A2(new_n227_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT25), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G183gat), .ZN(new_n240_));
  INV_X1    g039(.A(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT26), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G190gat), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n238_), .A2(new_n240_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n228_), .A2(new_n232_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT24), .A3(new_n234_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n221_), .A2(new_n223_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT24), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT92), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n254_), .A3(new_n251_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n248_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n218_), .B1(new_n236_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n252_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n245_), .A2(KEYINPUT83), .A3(new_n247_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT83), .B1(new_n245_), .B2(new_n247_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n224_), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n228_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT22), .B1(new_n228_), .B2(KEYINPUT84), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n232_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n262_), .A2(new_n265_), .A3(new_n234_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n209_), .A2(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n257_), .A2(KEYINPUT20), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n261_), .A2(new_n266_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n218_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n271_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n253_), .A2(new_n255_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n248_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n226_), .A2(new_n227_), .A3(new_n235_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n267_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n274_), .A2(KEYINPUT20), .A3(new_n275_), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n272_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT18), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT94), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G64gat), .B(G92gat), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n282_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  INV_X1    g094(.A(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n290_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n272_), .A2(new_n297_), .A3(new_n281_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n294_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n269_), .A2(new_n275_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n274_), .A2(KEYINPUT20), .A3(new_n271_), .A4(new_n280_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n293_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT98), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n293_), .A4(KEYINPUT98), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n298_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n299_), .B1(KEYINPUT27), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  OAI22_X1  g107(.A1(new_n308_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT3), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT2), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n308_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n311_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G141gat), .B(G148gat), .Z(new_n325_));
  NOR2_X1   g124(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(new_n321_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT1), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n324_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n331_));
  XOR2_X1   g130(.A(G22gat), .B(G50gat), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n331_), .A2(new_n332_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT89), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n334_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n331_), .A2(new_n332_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n340_), .B2(new_n333_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n330_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n344_), .B(new_n218_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n348_));
  OAI211_X1 g147(.A(G228gat), .B(G233gat), .C1(new_n348_), .C2(new_n267_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n343_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT91), .ZN(new_n351_));
  OAI22_X1  g150(.A1(new_n339_), .A2(new_n341_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n349_), .A3(new_n343_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n350_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(KEYINPUT91), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n356_), .B(new_n357_), .C1(new_n339_), .C2(new_n341_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  INV_X1    g159(.A(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(G15gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n362_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT85), .B(KEYINPUT30), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n261_), .A2(new_n266_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n367_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n372_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n370_), .A3(new_n366_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT86), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G134gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G127gat), .ZN(new_n380_));
  INV_X1    g179(.A(G113gat), .ZN(new_n381_));
  INV_X1    g180(.A(G120gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G127gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G134gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G113gat), .A2(G120gat), .ZN(new_n386_));
  AND4_X1   g185(.A1(new_n380_), .A2(new_n383_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n380_), .A2(new_n385_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT31), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n378_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n376_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G1gat), .B(G29gat), .Z(new_n395_));
  INV_X1    g194(.A(KEYINPUT0), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT0), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G57gat), .ZN(new_n401_));
  INV_X1    g200(.A(G57gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G85gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n401_), .A2(G85gat), .A3(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n389_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n330_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n324_), .A2(new_n329_), .A3(new_n389_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n324_), .A2(new_n389_), .A3(new_n329_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n389_), .B1(new_n324_), .B2(new_n329_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n330_), .A2(new_n416_), .A3(new_n409_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n412_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n408_), .B(new_n413_), .C1(new_n417_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT96), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n410_), .A2(new_n411_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n416_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n408_), .A4(new_n413_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n413_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n401_), .A2(G85gat), .A3(new_n403_), .ZN(new_n429_));
  AOI21_X1  g228(.A(G85gat), .B1(new_n401_), .B2(new_n403_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n422_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n394_), .A2(new_n433_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n307_), .A2(new_n359_), .A3(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n355_), .A2(new_n358_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n422_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n300_), .A2(new_n301_), .A3(new_n297_), .A4(KEYINPUT32), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n272_), .B(new_n281_), .C1(new_n293_), .C2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n437_), .A2(KEYINPUT97), .A3(new_n438_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n421_), .A2(KEYINPUT33), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n425_), .A2(new_n443_), .A3(new_n408_), .A4(new_n413_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n410_), .A2(new_n411_), .A3(new_n419_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n431_), .A2(KEYINPUT95), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT95), .B1(new_n431_), .B2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n418_), .A2(new_n412_), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n447_), .A2(new_n448_), .B1(new_n417_), .B2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n450_), .A3(new_n294_), .A4(new_n298_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n441_), .A2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n440_), .A2(new_n438_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT97), .B1(new_n453_), .B2(new_n437_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n436_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n437_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n282_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n457_), .A2(new_n297_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n295_), .B1(new_n458_), .B2(new_n305_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n456_), .B1(new_n459_), .B2(new_n299_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n394_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n435_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n464_));
  AND2_X1   g263(.A1(G230gat), .A2(G233gat), .ZN(new_n465_));
  AND3_X1   g264(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI22_X1  g267(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT64), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI221_X1 g270(.A(KEYINPUT64), .B1(KEYINPUT65), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AND2_X1   g272(.A1(G85gat), .A2(G92gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT8), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n479_), .A3(new_n476_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  AOI211_X1 g282(.A(new_n467_), .B(new_n466_), .C1(new_n483_), .C2(new_n474_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(KEYINPUT9), .ZN(new_n485_));
  OR2_X1    g284(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n486_));
  INV_X1    g285(.A(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n481_), .A2(new_n482_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G71gat), .B(G78gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(KEYINPUT11), .B2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n493_), .A3(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n491_), .A2(new_n492_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n484_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n473_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n479_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n497_), .A2(new_n498_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT67), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n491_), .A2(new_n499_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n465_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT68), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n501_), .B(new_n511_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n497_), .A2(KEYINPUT12), .A3(new_n498_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT12), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n465_), .B1(new_n491_), .B2(new_n499_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n509_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G120gat), .B(G148gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT5), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G176gat), .B(G204gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n509_), .A2(new_n519_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n524_), .B(KEYINPUT69), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(KEYINPUT13), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT13), .B1(new_n525_), .B2(new_n528_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n464_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(KEYINPUT70), .A3(new_n529_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT81), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT82), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G29gat), .B(G36gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT15), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT77), .B(G15gat), .Z(new_n548_));
  INV_X1    g347(.A(G22gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT77), .B(G15gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(G22gat), .ZN(new_n552_));
  INV_X1    g351(.A(G1gat), .ZN(new_n553_));
  INV_X1    g352(.A(G8gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G1gat), .B(G8gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n546_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT80), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT80), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n558_), .A2(new_n563_), .A3(new_n546_), .A4(new_n559_), .ZN(new_n564_));
  AOI221_X4 g363(.A(new_n543_), .B1(new_n547_), .B2(new_n560_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n561_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n542_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n541_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(new_n547_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n542_), .A3(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n562_), .A2(new_n564_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n571_), .B(KEYINPUT82), .C1(new_n572_), .C2(new_n542_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n540_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n540_), .A3(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n532_), .A2(new_n534_), .A3(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n463_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n510_), .A2(new_n512_), .A3(new_n547_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT35), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n491_), .B2(new_n546_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(KEYINPUT35), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n581_), .A2(KEYINPUT71), .A3(new_n585_), .A4(new_n588_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT36), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n592_), .A2(new_n593_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT73), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n599_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  AOI211_X1 g404(.A(KEYINPUT74), .B(new_n603_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n580_), .B(new_n598_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT76), .ZN(new_n608_));
  INV_X1    g407(.A(new_n591_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n589_), .B(new_n609_), .C1(new_n581_), .C2(new_n585_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n593_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n604_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT74), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n600_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(new_n580_), .A4(new_n598_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n597_), .B(KEYINPUT75), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n592_), .A2(new_n593_), .A3(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT37), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n608_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT16), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT78), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n560_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n499_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n628_), .B1(new_n631_), .B2(KEYINPUT79), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n632_), .B(KEYINPUT17), .C1(new_n628_), .C2(new_n631_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n634_), .B(new_n628_), .C1(new_n631_), .C2(KEYINPUT79), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n622_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n579_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n553_), .A3(new_n437_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n615_), .A2(new_n598_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n463_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n578_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n636_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n433_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n306_), .A2(KEYINPUT27), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n294_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n649_), .B(G8gat), .C1(new_n646_), .C2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT99), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT99), .ZN(new_n655_));
  INV_X1    g454(.A(new_n646_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n554_), .B1(new_n656_), .B2(new_n307_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n654_), .B(new_n655_), .C1(new_n649_), .C2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n638_), .A2(new_n554_), .A3(new_n307_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(KEYINPUT40), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n646_), .B2(new_n462_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n638_), .A2(new_n364_), .A3(new_n394_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1326gat));
  OAI21_X1  g468(.A(G22gat), .B1(new_n646_), .B2(new_n436_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT42), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n638_), .A2(new_n549_), .A3(new_n359_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n645_), .A2(new_n641_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n579_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n437_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n608_), .A2(new_n617_), .A3(new_n621_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n463_), .B2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n652_), .A2(new_n433_), .A3(new_n394_), .A4(new_n436_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT97), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n440_), .A2(new_n438_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n433_), .B2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n441_), .A3(new_n451_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n685_), .A2(new_n436_), .B1(new_n652_), .B2(new_n456_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n686_), .B2(new_n394_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n622_), .A3(new_n688_), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n578_), .B(new_n645_), .C1(new_n680_), .C2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n678_), .B1(new_n690_), .B2(KEYINPUT44), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n680_), .A2(new_n689_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n644_), .A3(new_n636_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT101), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n644_), .A4(new_n636_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n697_), .A2(G29gat), .A3(new_n437_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n677_), .B1(new_n696_), .B2(new_n698_), .ZN(G1328gat));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  INV_X1    g500(.A(new_n697_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n703_), .B2(new_n307_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n675_), .A2(G36gat), .A3(new_n652_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n700_), .B1(new_n704_), .B2(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n690_), .A2(new_n678_), .A3(KEYINPUT44), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT101), .B1(new_n693_), .B2(new_n694_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n307_), .B(new_n697_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT46), .A3(new_n707_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n709_), .A2(new_n714_), .ZN(G1329gat));
  NAND4_X1  g514(.A1(new_n696_), .A2(G43gat), .A3(new_n394_), .A4(new_n697_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n361_), .B1(new_n675_), .B2(new_n462_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n720_), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n676_), .A2(new_n723_), .A3(new_n359_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n697_), .A2(new_n359_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n723_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n726_), .A2(KEYINPUT103), .A3(new_n723_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n724_), .B1(new_n729_), .B2(new_n730_), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n532_), .A2(new_n534_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n637_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n637_), .A2(KEYINPUT104), .A3(new_n732_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n463_), .B2(new_n577_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738_));
  INV_X1    g537(.A(new_n577_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n687_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n735_), .A2(new_n736_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n735_), .A2(KEYINPUT106), .A3(new_n736_), .A4(new_n741_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n437_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n402_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n732_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(new_n577_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n750_));
  OR3_X1    g549(.A1(new_n750_), .A2(new_n402_), .A3(new_n433_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n747_), .A2(KEYINPUT107), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1332gat));
  OAI21_X1  g555(.A(G64gat), .B1(new_n750_), .B2(new_n652_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n744_), .A2(new_n745_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n652_), .A2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g562(.A(G71gat), .B1(new_n750_), .B2(new_n462_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT49), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n462_), .A2(G71gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n760_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1334gat));
  OAI21_X1  g568(.A(G78gat), .B1(new_n750_), .B2(new_n436_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n436_), .A2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n760_), .B2(new_n773_), .ZN(G1335gat));
  NAND3_X1  g573(.A1(new_n692_), .A2(new_n636_), .A3(new_n749_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n433_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n674_), .A2(new_n732_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n405_), .A3(new_n437_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n775_), .B2(new_n652_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n778_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n652_), .A2(G92gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT112), .Z(G1337gat));
  INV_X1    g584(.A(new_n777_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n394_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n741_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n778_), .A2(KEYINPUT113), .A3(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  OAI21_X1  g592(.A(G99gat), .B1(new_n775_), .B2(new_n462_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT115), .B(KEYINPUT51), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n794_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT114), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n798_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  INV_X1    g602(.A(new_n799_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n798_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n797_), .B1(new_n802_), .B2(new_n805_), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n778_), .A2(new_n487_), .A3(new_n359_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  INV_X1    g607(.A(new_n775_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n359_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(G106gat), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT52), .B(new_n487_), .C1(new_n809_), .C2(new_n359_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n807_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT53), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n807_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1339gat));
  NOR3_X1   g616(.A1(new_n577_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n679_), .A2(new_n818_), .A3(new_n645_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n525_), .A2(new_n528_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n572_), .A2(new_n543_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n566_), .A2(new_n543_), .A3(new_n570_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n537_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n538_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n569_), .A2(new_n540_), .A3(new_n573_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n525_), .B1(new_n831_), .B2(new_n574_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n527_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n515_), .A2(new_n506_), .A3(new_n500_), .A4(new_n517_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n465_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n515_), .A2(KEYINPUT55), .A3(new_n517_), .A4(new_n518_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n519_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n836_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT116), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n465_), .A2(new_n834_), .B1(new_n519_), .B2(new_n837_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n836_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n833_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(KEYINPUT117), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n832_), .B1(new_n845_), .B2(KEYINPUT56), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(KEYINPUT117), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n830_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n822_), .B1(new_n849_), .B2(new_n642_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n842_), .B1(new_n841_), .B2(new_n836_), .ZN(new_n851_));
  AND4_X1   g650(.A1(new_n842_), .A2(new_n835_), .A3(new_n836_), .A4(new_n838_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n527_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(KEYINPUT56), .ZN(new_n855_));
  INV_X1    g654(.A(new_n525_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n829_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(KEYINPUT57), .A3(new_n641_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n853_), .A2(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n844_), .A2(new_n847_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n828_), .A2(new_n525_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n861_), .A2(new_n862_), .A3(KEYINPUT58), .A4(new_n863_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n622_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n850_), .A2(new_n860_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n821_), .B1(new_n869_), .B2(new_n636_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n307_), .A2(new_n359_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n437_), .A3(new_n394_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n381_), .A3(new_n577_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n872_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n622_), .A2(new_n867_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n642_), .B1(new_n858_), .B2(new_n829_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n878_), .A2(new_n866_), .B1(new_n879_), .B2(KEYINPUT57), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n645_), .B1(new_n880_), .B2(new_n850_), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT59), .B(new_n877_), .C1(new_n881_), .C2(new_n821_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n739_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n874_), .B1(new_n883_), .B2(new_n381_), .ZN(G1340gat));
  AOI21_X1  g683(.A(new_n748_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n860_), .A2(new_n868_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n879_), .A2(KEYINPUT57), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n636_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n821_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n877_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n748_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n893_));
  OAI22_X1  g692(.A1(new_n885_), .A2(new_n382_), .B1(new_n891_), .B2(new_n893_), .ZN(G1341gat));
  NAND3_X1  g693(.A1(new_n873_), .A2(new_n384_), .A3(new_n645_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n636_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n384_), .ZN(G1342gat));
  NOR2_X1   g696(.A1(new_n679_), .A2(new_n379_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n882_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT59), .B1(new_n890_), .B2(new_n877_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n379_), .B1(new_n891_), .B2(new_n641_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n898_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G134gat), .B1(new_n873_), .B2(new_n642_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT118), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n908_), .ZN(G1343gat));
  NOR2_X1   g708(.A1(new_n436_), .A2(new_n394_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n911_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n307_), .A2(new_n433_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n577_), .A3(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n732_), .A3(new_n913_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g716(.A1(new_n890_), .A2(new_n645_), .A3(new_n910_), .A4(new_n913_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT119), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n912_), .A2(new_n920_), .A3(new_n645_), .A4(new_n913_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT61), .B(G155gat), .Z(new_n922_));
  AND3_X1   g721(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1346gat));
  NAND2_X1  g724(.A1(new_n912_), .A2(new_n913_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G162gat), .B1(new_n926_), .B2(new_n679_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n642_), .A2(new_n320_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1347gat));
  AOI21_X1  g728(.A(new_n359_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n652_), .A2(new_n434_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n739_), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n930_), .A2(new_n229_), .A3(new_n231_), .A4(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n933_), .B(KEYINPUT120), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n930_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n935_), .B1(new_n938_), .B2(G169gat), .ZN(new_n939_));
  AOI211_X1 g738(.A(KEYINPUT62), .B(new_n228_), .C1(new_n930_), .C2(new_n937_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n934_), .B1(new_n939_), .B2(new_n940_), .ZN(G1348gat));
  NAND2_X1  g740(.A1(new_n930_), .A2(new_n931_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n748_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n943_), .A2(new_n944_), .A3(new_n232_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT121), .B(G176gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n943_), .B2(new_n946_), .ZN(G1349gat));
  AND2_X1   g746(.A1(new_n238_), .A2(new_n240_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n930_), .A2(new_n948_), .A3(new_n645_), .A4(new_n931_), .ZN(new_n949_));
  NOR4_X1   g748(.A1(new_n870_), .A2(new_n359_), .A3(new_n636_), .A4(new_n932_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n237_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(KEYINPUT122), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n953_), .B(new_n949_), .C1(new_n950_), .C2(new_n237_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n954_), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n942_), .B2(new_n679_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n642_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n942_), .B2(new_n957_), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n652_), .A2(new_n437_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n912_), .A2(new_n577_), .A3(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n961_));
  INV_X1    g760(.A(G197gat), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n960_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n961_), .B1(new_n960_), .B2(new_n962_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n960_), .A2(new_n962_), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n963_), .A2(new_n964_), .A3(new_n965_), .ZN(G1352gat));
  AND3_X1   g765(.A1(new_n890_), .A2(new_n910_), .A3(new_n959_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(new_n732_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g768(.A(KEYINPUT125), .ZN(new_n970_));
  NOR2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  INV_X1    g770(.A(new_n971_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n636_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(KEYINPUT124), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n967_), .A2(new_n970_), .A3(new_n972_), .A4(new_n974_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n912_), .A2(new_n959_), .A3(new_n974_), .ZN(new_n976_));
  OAI21_X1  g775(.A(KEYINPUT125), .B1(new_n976_), .B2(new_n971_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n971_), .ZN(new_n978_));
  AND3_X1   g777(.A1(new_n975_), .A2(new_n977_), .A3(new_n978_), .ZN(G1354gat));
  NAND2_X1  g778(.A1(new_n967_), .A2(new_n642_), .ZN(new_n980_));
  XOR2_X1   g779(.A(KEYINPUT126), .B(G218gat), .Z(new_n981_));
  NOR2_X1   g780(.A1(new_n679_), .A2(new_n981_), .ZN(new_n982_));
  AOI22_X1  g781(.A1(new_n980_), .A2(new_n981_), .B1(new_n967_), .B2(new_n982_), .ZN(G1355gat));
endmodule


