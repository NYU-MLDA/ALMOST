//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT93), .Z(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT90), .B1(new_n205_), .B2(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT90), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT21), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT92), .Z(new_n214_));
  OR2_X1    g013(.A1(new_n211_), .A2(KEYINPUT21), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT91), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n208_), .A2(G204gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n210_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n212_), .B1(KEYINPUT21), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n214_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT23), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT94), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT95), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n232_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n227_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G169gat), .ZN(new_n238_));
  INV_X1    g037(.A(G176gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n240_), .A2(new_n233_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT96), .Z(new_n242_));
  OAI21_X1  g041(.A(new_n226_), .B1(G183gat), .B2(G190gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT97), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n221_), .B1(new_n237_), .B2(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n215_), .A2(new_n216_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n215_), .A2(new_n216_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n220_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n213_), .B(KEYINPUT92), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(new_n243_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n227_), .A2(new_n234_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n230_), .A2(KEYINPUT84), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT84), .B1(new_n255_), .B2(G190gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(new_n228_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n252_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT20), .B1(new_n251_), .B2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n204_), .B1(new_n246_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n221_), .A2(new_n237_), .A3(new_n245_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n203_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n261_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT18), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(G64gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(G92gat), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n270_), .A3(new_n265_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n272_), .A2(KEYINPUT98), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT98), .B1(new_n272_), .B2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G127gat), .B(G134gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT86), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT87), .Z(new_n281_));
  NOR2_X1   g080(.A1(new_n277_), .A2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G141gat), .A2(G148gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G155gat), .B(G162gat), .Z(new_n288_));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT88), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n284_), .B(KEYINPUT3), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n286_), .B(KEYINPUT2), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n288_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n280_), .B(KEYINPUT87), .ZN(new_n300_));
  INV_X1    g099(.A(new_n282_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n283_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n292_), .A2(new_n293_), .B1(new_n297_), .B2(new_n288_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n279_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT4), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n303_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G57gat), .B(G85gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G29gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT33), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n315_), .A2(KEYINPUT33), .A3(new_n320_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n320_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n303_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n308_), .A2(new_n312_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n325_), .B(new_n326_), .C1(new_n327_), .C2(new_n310_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n313_), .A2(new_n325_), .A3(new_n314_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(KEYINPUT100), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT100), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n315_), .A2(new_n332_), .A3(new_n320_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(new_n246_), .A2(new_n204_), .A3(new_n259_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n264_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(KEYINPUT32), .A3(new_n270_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n266_), .ZN(new_n341_));
  OAI22_X1  g140(.A1(new_n276_), .A2(new_n329_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT28), .B1(new_n299_), .B2(KEYINPUT29), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n304_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT89), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n349_), .A3(new_n346_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G228gat), .ZN(new_n354_));
  INV_X1    g153(.A(G233gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n299_), .A2(KEYINPUT29), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n251_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n357_), .A3(new_n251_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G22gat), .B(G50gat), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n361_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n362_), .B1(new_n365_), .B2(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n352_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n348_), .A2(new_n350_), .A3(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n353_), .A2(new_n364_), .A3(new_n366_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n364_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n348_), .A2(new_n350_), .A3(new_n367_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  INV_X1    g174(.A(new_n273_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n270_), .B1(new_n260_), .B2(new_n265_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT102), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT102), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n380_), .B(new_n375_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT101), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n338_), .A2(new_n382_), .A3(new_n271_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n246_), .A2(new_n259_), .A3(new_n204_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n271_), .B1(new_n384_), .B2(new_n336_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT101), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n376_), .A2(new_n375_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n379_), .A2(new_n381_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n374_), .B1(new_n333_), .B2(new_n331_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n342_), .A2(new_n374_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n283_), .A2(new_n302_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G71gat), .B(G99gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(G15gat), .B(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n392_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n258_), .B(KEYINPUT30), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n400_), .A2(new_n401_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n403_), .A2(KEYINPUT31), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT31), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n258_), .B(KEYINPUT30), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT85), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n408_), .B2(new_n402_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n399_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT31), .B1(new_n403_), .B2(new_n404_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(new_n402_), .A3(new_n406_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n398_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n369_), .A2(new_n373_), .A3(new_n410_), .A4(new_n413_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n333_), .B2(new_n331_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT103), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n389_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n389_), .B2(new_n417_), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n391_), .A2(new_n415_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G85gat), .B(G92gat), .Z(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT9), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G99gat), .A2(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT65), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT6), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n425_), .ZN(new_n431_));
  OAI221_X1 g230(.A(new_n423_), .B1(KEYINPUT9), .B2(new_n424_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT10), .B(G99gat), .Z(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n433_), .A2(KEYINPUT64), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT64), .B1(new_n433_), .B2(new_n434_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n431_), .A2(new_n430_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT66), .A2(G99gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n434_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT7), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n444_), .A3(new_n434_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n439_), .B(new_n422_), .C1(new_n440_), .C2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT6), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n426_), .A2(KEYINPUT67), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n425_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n425_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n426_), .A2(KEYINPUT67), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(KEYINPUT6), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n451_), .A2(new_n443_), .A3(new_n445_), .A4(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n439_), .B1(new_n456_), .B2(new_n422_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n447_), .B1(new_n457_), .B2(KEYINPUT68), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n459_), .B(new_n439_), .C1(new_n456_), .C2(new_n422_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n438_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT69), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n467_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n468_), .A2(KEYINPUT15), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT15), .B1(new_n468_), .B2(new_n469_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n438_), .B(KEYINPUT69), .C1(new_n458_), .C2(new_n460_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n463_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G232gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT34), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT35), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(KEYINPUT35), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n432_), .A2(new_n437_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n422_), .A2(new_n439_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n431_), .A2(new_n430_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n446_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n456_), .A2(new_n422_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT8), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n485_), .B2(new_n459_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n460_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n479_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n468_), .A2(new_n469_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n474_), .A2(new_n477_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n477_), .B1(new_n474_), .B2(new_n490_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT79), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G134gat), .B(G162gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT78), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G190gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G218gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n498_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n493_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  OAI221_X1 g302(.A(KEYINPUT79), .B1(new_n503_), .B2(new_n499_), .C1(new_n491_), .C2(new_n492_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n502_), .A2(KEYINPUT105), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT105), .B1(new_n502_), .B2(new_n504_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT106), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT106), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G15gat), .B(G22gat), .Z(new_n511_));
  NAND2_X1  g310(.A1(G1gat), .A2(G8gat), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(KEYINPUT14), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT81), .ZN(new_n514_));
  XOR2_X1   g313(.A(G1gat), .B(G8gat), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n513_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G231gat), .A2(G233gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G71gat), .B(G78gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(KEYINPUT11), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n526_), .A3(KEYINPUT11), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n523_), .B(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G183gat), .B(G211gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(G127gat), .B(G155gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n537_), .B(KEYINPUT17), .Z(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(KEYINPUT70), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n529_), .A2(new_n530_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n523_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n523_), .A2(new_n544_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n545_), .A2(KEYINPUT17), .A3(new_n537_), .A4(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n539_), .A2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n421_), .A2(new_n510_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n463_), .A2(new_n473_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n461_), .A2(new_n531_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n550_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n438_), .B(new_n541_), .C1(new_n458_), .C2(new_n460_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n555_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n556_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n552_), .A2(new_n554_), .A3(KEYINPUT71), .A4(new_n557_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G120gat), .B(G148gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT72), .B(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT5), .B(G176gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  NAND4_X1  g368(.A1(new_n560_), .A2(new_n563_), .A3(new_n564_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT73), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n560_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n573_));
  INV_X1    g372(.A(new_n569_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n573_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n571_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT74), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n570_), .A2(KEYINPUT73), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n577_), .A2(new_n582_), .A3(new_n584_), .A4(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n472_), .A2(new_n521_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n516_), .A2(new_n520_), .A3(new_n489_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n489_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n521_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n592_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n598_), .B2(new_n593_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(G169gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n208_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(KEYINPUT83), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n599_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n590_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n549_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT107), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT107), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n549_), .A2(new_n610_), .A3(new_n607_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n334_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G1gat), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n421_), .A2(new_n605_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n588_), .A2(new_n589_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT80), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n502_), .A2(new_n619_), .A3(new_n504_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n618_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n502_), .A2(new_n504_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT80), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n502_), .A2(new_n619_), .A3(new_n504_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(KEYINPUT37), .A3(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n622_), .A2(new_n626_), .A3(new_n548_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n616_), .A2(new_n617_), .A3(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n334_), .A2(G1gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n615_), .A2(new_n631_), .A3(new_n632_), .ZN(G1324gat));
  OR3_X1    g432(.A1(new_n628_), .A2(G8gat), .A3(new_n389_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G8gat), .B1(new_n608_), .B2(new_n389_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(KEYINPUT39), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(KEYINPUT39), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g438(.A1(new_n628_), .A2(G15gat), .A3(new_n414_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n612_), .A2(new_n415_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n641_), .B2(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  OR3_X1    g443(.A1(new_n628_), .A2(G22gat), .A3(new_n374_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n374_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n609_), .A2(new_n611_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G22gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT108), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n650_), .A3(G22gat), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n649_), .A2(KEYINPUT42), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT42), .B1(new_n649_), .B2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n645_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n507_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n548_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n616_), .A2(new_n617_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n613_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n622_), .A2(new_n626_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n421_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT110), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT110), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n421_), .A2(new_n664_), .A3(new_n660_), .A4(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n421_), .A2(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n590_), .A2(new_n606_), .A3(new_n548_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT109), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n670_), .A3(KEYINPUT44), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(G29gat), .A3(new_n613_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n670_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n659_), .B1(new_n672_), .B2(new_n674_), .ZN(G1328gat));
  INV_X1    g474(.A(new_n389_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G36gat), .B1(new_n677_), .B2(new_n673_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n389_), .A2(G36gat), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n657_), .A2(KEYINPUT111), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT111), .B1(new_n657_), .B2(new_n679_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n678_), .A2(new_n685_), .A3(KEYINPUT46), .A4(new_n682_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  NAND3_X1  g489(.A1(new_n671_), .A2(G43gat), .A3(new_n415_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n657_), .A2(new_n414_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n691_), .A2(new_n673_), .B1(G43gat), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1330gat));
  AOI21_X1  g494(.A(G50gat), .B1(new_n658_), .B2(new_n646_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n671_), .A2(G50gat), .A3(new_n646_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n674_), .ZN(G1331gat));
  AND2_X1   g497(.A1(new_n421_), .A2(new_n606_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n590_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n627_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n613_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n510_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n548_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n700_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n613_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n708_), .B2(new_n703_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n707_), .B2(new_n676_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT48), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n676_), .A2(new_n710_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT113), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n702_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n707_), .B2(new_n415_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT49), .Z(new_n719_));
  NAND3_X1  g518(.A1(new_n702_), .A2(new_n717_), .A3(new_n415_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1334gat));
  INV_X1    g520(.A(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n707_), .B2(new_n646_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n702_), .A2(new_n722_), .A3(new_n646_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1335gat));
  NAND3_X1  g525(.A1(new_n590_), .A2(new_n606_), .A3(new_n706_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT114), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n668_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n334_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n656_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n700_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(G85gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n733_), .A3(new_n613_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1336gat));
  NAND2_X1  g534(.A1(new_n676_), .A2(G92gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT115), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n729_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G92gat), .B1(new_n732_), .B2(new_n676_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1337gat));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n668_), .A2(new_n415_), .A3(new_n728_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G99gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n415_), .A2(new_n433_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n700_), .A2(new_n731_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n741_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n746_), .A3(new_n741_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT116), .B(new_n745_), .C1(new_n742_), .C2(G99gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n747_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n750_), .A2(new_n753_), .ZN(G1338gat));
  OAI21_X1  g553(.A(G106gat), .B1(new_n729_), .B2(new_n374_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n374_), .A2(G106gat), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n699_), .A2(new_n590_), .A3(new_n656_), .A4(new_n758_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT117), .Z(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT52), .B(G106gat), .C1(new_n729_), .C2(new_n374_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n757_), .A2(new_n760_), .A3(new_n764_), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  NOR3_X1   g565(.A1(new_n676_), .A2(new_n334_), .A3(new_n416_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(KEYINPUT124), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(KEYINPUT124), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(KEYINPUT59), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n599_), .A2(new_n603_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n593_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n591_), .A2(new_n592_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n603_), .B1(new_n598_), .B2(new_n773_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(KEYINPUT119), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n603_), .C1(new_n598_), .C2(new_n773_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n772_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n570_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n560_), .A2(new_n781_), .A3(new_n564_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n552_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n552_), .A2(new_n555_), .A3(new_n554_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n783_), .A2(KEYINPUT55), .B1(new_n784_), .B2(new_n562_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n569_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n788_), .B(new_n569_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n780_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT121), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT58), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  OAI221_X1 g592(.A(new_n780_), .B1(new_n791_), .B2(KEYINPUT58), .C1(new_n787_), .C2(new_n789_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n661_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n577_), .A2(new_n582_), .A3(new_n779_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n782_), .A2(new_n785_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n797_), .B(KEYINPUT56), .C1(new_n798_), .C2(new_n569_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n788_), .B1(new_n786_), .B2(KEYINPUT118), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n605_), .A2(new_n570_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n507_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n803_), .A2(KEYINPUT122), .A3(new_n805_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n795_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n655_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT120), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n507_), .B1(new_n796_), .B2(new_n802_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n804_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n548_), .B1(new_n810_), .B2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n627_), .A2(new_n606_), .A3(new_n589_), .A4(new_n588_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT54), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n617_), .A2(new_n820_), .A3(new_n606_), .A4(new_n627_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n771_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT125), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n661_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n809_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT122), .B1(new_n803_), .B2(new_n805_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n804_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT120), .B(new_n507_), .C1(new_n796_), .C2(new_n802_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n706_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n819_), .A2(new_n821_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n771_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n824_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n767_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n605_), .A2(G113gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT126), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n768_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n605_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n844_), .A2(KEYINPUT123), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(KEYINPUT123), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n840_), .A2(new_n842_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT60), .B1(new_n590_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(KEYINPUT60), .B2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n843_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n590_), .B1(new_n843_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n824_), .B2(new_n836_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT127), .B(new_n851_), .C1(new_n854_), .C2(new_n848_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT127), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n617_), .B1(new_n838_), .B2(KEYINPUT59), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n848_), .B1(new_n837_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n851_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n855_), .A2(new_n860_), .ZN(G1341gat));
  NAND3_X1  g660(.A1(new_n837_), .A2(new_n548_), .A3(new_n839_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G127gat), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n706_), .A2(G127gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n838_), .B2(new_n864_), .ZN(G1342gat));
  NAND3_X1  g664(.A1(new_n837_), .A2(new_n661_), .A3(new_n839_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G134gat), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n510_), .A2(G134gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n838_), .B2(new_n868_), .ZN(G1343gat));
  NOR4_X1   g668(.A1(new_n676_), .A2(new_n334_), .A3(new_n374_), .A4(new_n415_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n834_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n605_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n590_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n706_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  INV_X1    g678(.A(new_n661_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G162gat), .B1(new_n871_), .B2(new_n880_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n510_), .A2(G162gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n871_), .B2(new_n882_), .ZN(G1347gat));
  NOR3_X1   g682(.A1(new_n389_), .A2(new_n613_), .A3(new_n416_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n834_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n605_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G169gat), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n238_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n890_), .B(new_n891_), .C1(new_n892_), .C2(new_n887_), .ZN(G1348gat));
  NOR2_X1   g692(.A1(new_n885_), .A2(new_n617_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n239_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n885_), .A2(new_n706_), .ZN(new_n896_));
  MUX2_X1   g695(.A(G183gat), .B(new_n229_), .S(new_n896_), .Z(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n885_), .B2(new_n880_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n705_), .A2(new_n230_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n885_), .B2(new_n899_), .ZN(G1351gat));
  NOR4_X1   g699(.A1(new_n389_), .A2(new_n613_), .A3(new_n374_), .A4(new_n415_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n834_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n606_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n208_), .ZN(G1352gat));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n617_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n205_), .ZN(G1353gat));
  NAND3_X1  g705(.A1(new_n834_), .A2(new_n548_), .A3(new_n901_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  AND2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n907_), .B2(new_n908_), .ZN(G1354gat));
  OAI21_X1  g710(.A(G218gat), .B1(new_n902_), .B2(new_n880_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n510_), .A2(G218gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n902_), .B2(new_n913_), .ZN(G1355gat));
endmodule


