//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  AND2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n205_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G141gat), .B(G148gat), .Z(new_n213_));
  INV_X1    g012(.A(KEYINPUT85), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(new_n204_), .B2(KEYINPUT1), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n203_), .A3(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n204_), .A2(new_n214_), .A3(KEYINPUT1), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n213_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G22gat), .B(G50gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n219_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n222_), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT91), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT91), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n228_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G197gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT87), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G197gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G204gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G197gat), .A2(G204gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n249_));
  INV_X1    g048(.A(G204gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n239_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n236_), .B1(G197gat), .B2(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n235_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n246_), .B1(new_n249_), .B2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n220_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(G228gat), .A3(G233gat), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n226_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(KEYINPUT89), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT89), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(new_n246_), .C1(new_n249_), .C2(new_n254_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n259_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n258_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n231_), .B(new_n234_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT91), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n258_), .A2(new_n263_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n264_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n258_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n269_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G71gat), .B(G99gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT25), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G183gat), .ZN(new_n280_));
  INV_X1    g079(.A(G183gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT25), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n282_), .A3(KEYINPUT78), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n281_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT26), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT26), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n289_), .A3(KEYINPUT79), .ZN(new_n290_));
  OR3_X1    g089(.A1(new_n288_), .A2(KEYINPUT79), .A3(KEYINPUT26), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n285_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n293_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT23), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  INV_X1    g097(.A(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT81), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n300_), .A2(new_n302_), .A3(KEYINPUT24), .A4(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n300_), .A2(new_n302_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n297_), .B(new_n304_), .C1(new_n305_), .C2(KEYINPUT24), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n294_), .A2(new_n295_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n297_), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n303_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n299_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n307_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n285_), .A2(new_n292_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT80), .ZN(new_n317_));
  INV_X1    g116(.A(new_n306_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n285_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT30), .B1(new_n320_), .B2(new_n313_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n278_), .B1(new_n315_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n313_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n308_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n295_), .A2(new_n306_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n314_), .B1(new_n325_), .B2(new_n319_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT30), .ZN(new_n327_));
  INV_X1    g126(.A(new_n278_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n322_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n330_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n275_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n328_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n315_), .A2(new_n321_), .A3(new_n278_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n322_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(KEYINPUT83), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G134gat), .Z(new_n340_));
  INV_X1    g139(.A(G120gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G113gat), .ZN(new_n342_));
  INV_X1    g141(.A(G113gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G120gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n333_), .A2(new_n339_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n337_), .A2(new_n338_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n275_), .A3(new_n351_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT0), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G57gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(G57gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n358_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n360_), .A2(G57gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G85gat), .A3(new_n361_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n349_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n226_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n372_), .B2(KEYINPUT4), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n212_), .A2(new_n219_), .A3(new_n349_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(KEYINPUT95), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT95), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n226_), .A2(new_n376_), .A3(new_n371_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n378_), .B2(KEYINPUT4), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n370_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n368_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n369_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n382_), .B(new_n367_), .C1(new_n384_), .C2(new_n373_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n354_), .A2(new_n357_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n287_), .A2(new_n289_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT92), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n287_), .A2(new_n289_), .A3(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n280_), .A2(new_n282_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n397_), .A2(new_n297_), .A3(new_n304_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT93), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n312_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n298_), .A2(KEYINPUT22), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G169gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n405_), .A3(new_n299_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n303_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT93), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n402_), .A2(new_n408_), .A3(new_n309_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n400_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT20), .B1(new_n410_), .B2(new_n255_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n260_), .B(new_n262_), .C1(new_n307_), .C2(new_n314_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n412_), .B2(KEYINPUT94), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n323_), .A2(new_n414_), .A3(new_n260_), .A4(new_n262_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n391_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n260_), .A2(new_n262_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n326_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT20), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n419_), .B1(new_n410_), .B2(new_n255_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n391_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G64gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G92gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n416_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT94), .B1(new_n417_), .B2(new_n326_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n411_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n415_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n391_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n426_), .B1(new_n433_), .B2(new_n421_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n389_), .B1(new_n428_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n416_), .B2(new_n422_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n418_), .A2(new_n420_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n432_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n438_), .B(new_n426_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(KEYINPUT27), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT99), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT99), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n443_), .A3(new_n440_), .ZN(new_n444_));
  AND4_X1   g243(.A1(new_n274_), .A2(new_n387_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n353_), .A2(KEYINPUT84), .A3(new_n356_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT84), .B1(new_n353_), .B2(new_n356_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n274_), .A2(new_n386_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n435_), .A2(new_n449_), .A3(new_n440_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n274_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n433_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n385_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n374_), .A2(KEYINPUT95), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n349_), .B1(new_n212_), .B2(new_n219_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n377_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT4), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n373_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n380_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n368_), .A2(new_n453_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n370_), .B1(new_n456_), .B2(new_n383_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n459_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n367_), .B1(new_n378_), .B2(new_n370_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n461_), .A2(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n436_), .A2(new_n452_), .A3(new_n454_), .A4(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n426_), .A2(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n438_), .B(new_n469_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n422_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n386_), .B(new_n470_), .C1(new_n471_), .C2(new_n469_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n451_), .B1(new_n467_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n450_), .B1(new_n473_), .B2(KEYINPUT96), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n475_));
  AOI211_X1 g274(.A(new_n475_), .B(new_n451_), .C1(new_n467_), .C2(new_n472_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n448_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT98), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT98), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n448_), .B(new_n479_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n445_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G85gat), .B(G92gat), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(KEYINPUT9), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT64), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT10), .B(G99gat), .Z(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT6), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(new_n490_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT7), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n483_), .A2(new_n499_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n486_), .A2(new_n492_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n491_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT65), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n496_), .A2(new_n504_), .A3(new_n491_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n483_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n499_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G29gat), .B(G36gat), .Z(new_n510_));
  XOR2_X1   g309(.A(G43gat), .B(G50gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT15), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n501_), .A2(new_n512_), .A3(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT69), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n514_), .A2(new_n515_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT70), .ZN(new_n527_));
  INV_X1    g326(.A(G134gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G162gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n522_), .A2(new_n524_), .B1(new_n525_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n531_), .B(new_n525_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n524_), .A3(new_n522_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n481_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G176gat), .B(G204gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G71gat), .B(G78gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(KEYINPUT11), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n486_), .A2(new_n492_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n498_), .A2(new_n500_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n483_), .B1(new_n502_), .B2(KEYINPUT65), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT8), .B1(new_n552_), .B2(new_n505_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n548_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n548_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n501_), .A2(new_n508_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n554_), .A2(new_n556_), .B1(KEYINPUT67), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n509_), .A2(new_n548_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n558_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n559_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n543_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n554_), .A2(new_n556_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n562_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n559_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n565_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n542_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT13), .ZN(new_n574_));
  XOR2_X1   g373(.A(G15gat), .B(G22gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT72), .B(G1gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(G8gat), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n575_), .B1(new_n577_), .B2(KEYINPUT14), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n202_), .ZN(new_n579_));
  INV_X1    g378(.A(G8gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n578_), .A2(new_n202_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n202_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(G8gat), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n512_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n584_), .ZN(new_n587_));
  AOI21_X1  g386(.A(G8gat), .B1(new_n582_), .B2(new_n583_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n512_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT75), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n591_), .A3(new_n512_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n586_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT76), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT76), .ZN(new_n596_));
  INV_X1    g395(.A(new_n594_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n591_), .B1(new_n585_), .B2(new_n512_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n512_), .ZN(new_n599_));
  AOI211_X1 g398(.A(KEYINPUT75), .B(new_n599_), .C1(new_n581_), .C2(new_n584_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n596_), .B(new_n597_), .C1(new_n601_), .C2(new_n586_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n585_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n590_), .A2(new_n592_), .B1(new_n513_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n594_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n595_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(G141gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT77), .B(G113gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n595_), .A2(new_n602_), .A3(new_n605_), .A4(new_n610_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n574_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n585_), .B(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(new_n548_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n548_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(KEYINPUT74), .A3(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n620_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n618_), .A2(KEYINPUT74), .A3(new_n619_), .A4(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n618_), .A2(new_n619_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n626_), .A3(new_n625_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n615_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n537_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n202_), .B1(new_n636_), .B2(new_n386_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT101), .ZN(new_n638_));
  INV_X1    g437(.A(new_n614_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT71), .ZN(new_n640_));
  INV_X1    g439(.A(new_n535_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n640_), .B(KEYINPUT37), .C1(new_n641_), .C2(new_n532_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n640_), .A2(KEYINPUT37), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(KEYINPUT37), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n533_), .A2(new_n535_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n631_), .A2(new_n633_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n574_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n481_), .A2(new_n639_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n386_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n576_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT38), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT102), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n653_), .A2(new_n654_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT100), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n638_), .A2(new_n656_), .A3(new_n658_), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n442_), .A2(new_n444_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n650_), .A2(new_n580_), .A3(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n537_), .A2(new_n660_), .A3(new_n635_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n662_), .A2(new_n663_), .A3(G8gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n662_), .B2(G8gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT103), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n668_), .B(new_n661_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g470(.A(G15gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n448_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n636_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT41), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n650_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n636_), .B2(new_n451_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT42), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n650_), .A2(new_n678_), .A3(new_n451_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  NOR2_X1   g481(.A1(new_n615_), .A2(new_n647_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n481_), .B2(new_n646_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n481_), .A2(KEYINPUT43), .A3(new_n646_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(KEYINPUT104), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n481_), .A2(new_n687_), .A3(KEYINPUT43), .A4(new_n646_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n683_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(G29gat), .A3(new_n386_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  INV_X1    g490(.A(new_n646_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n478_), .A2(new_n480_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n691_), .B(new_n692_), .C1(new_n693_), .C2(new_n445_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n687_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n685_), .A2(KEYINPUT104), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n684_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n683_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n536_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n647_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT105), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(new_n574_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n481_), .A2(new_n639_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n651_), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n690_), .A2(new_n698_), .B1(G29gat), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT106), .ZN(G1328gat));
  NAND2_X1  g506(.A1(new_n689_), .A2(new_n660_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G36gat), .B1(new_n708_), .B2(new_n698_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n660_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n702_), .A2(new_n703_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT107), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n702_), .A2(new_n703_), .A3(new_n714_), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT45), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n709_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n709_), .A2(new_n717_), .A3(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  NOR2_X1   g521(.A1(new_n354_), .A2(new_n357_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n689_), .A2(G43gat), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n704_), .A2(new_n448_), .ZN(new_n725_));
  OAI22_X1  g524(.A1(new_n724_), .A2(new_n698_), .B1(G43gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g526(.A1(new_n704_), .A2(new_n274_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(G50gat), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n689_), .A2(G50gat), .A3(new_n451_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n698_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n574_), .A2(new_n614_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n481_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n648_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT108), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n386_), .ZN(new_n738_));
  INV_X1    g537(.A(G57gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NOR4_X1   g539(.A1(new_n481_), .A2(new_n536_), .A3(new_n634_), .A4(new_n734_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(G57gat), .A3(new_n386_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g544(.A(G64gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n741_), .B2(new_n660_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT48), .Z(new_n748_));
  NAND2_X1  g547(.A1(new_n660_), .A2(new_n746_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT111), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n737_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n741_), .B2(new_n673_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n737_), .A2(new_n753_), .A3(new_n673_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n741_), .B2(new_n451_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT50), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n737_), .A2(new_n759_), .A3(new_n451_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n734_), .A2(new_n647_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n697_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n651_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n735_), .A2(new_n701_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n358_), .A3(new_n386_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n710_), .ZN(new_n770_));
  INV_X1    g569(.A(G92gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(new_n771_), .A3(new_n660_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n765_), .B2(new_n448_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n767_), .A2(new_n723_), .A3(new_n487_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n488_), .A3(new_n451_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n451_), .B(new_n764_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n778_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  AOI21_X1  g586(.A(new_n610_), .B1(new_n604_), .B2(new_n597_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n597_), .B2(new_n593_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n613_), .A2(new_n789_), .A3(new_n572_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n560_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n564_), .B2(KEYINPUT55), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n568_), .A2(KEYINPUT55), .A3(new_n559_), .A4(new_n569_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT56), .B(new_n543_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n570_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n793_), .A3(new_n791_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n543_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n790_), .B1(new_n796_), .B2(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n802_));
  AOI21_X1  g601(.A(new_n646_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n790_), .B(KEYINPUT58), .C1(new_n796_), .C2(new_n800_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n799_), .A2(new_n543_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n795_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n790_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n803_), .A2(new_n806_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n795_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n799_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n543_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n809_), .A3(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n564_), .A2(new_n565_), .A3(new_n543_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n573_), .A2(new_n613_), .A3(new_n789_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n573_), .A2(new_n613_), .A3(new_n789_), .A4(KEYINPUT115), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n536_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n812_), .B1(new_n825_), .B2(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n823_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n536_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n634_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n614_), .B1(KEYINPUT113), .B2(KEYINPUT54), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n649_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n832_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n648_), .A2(new_n574_), .A3(new_n833_), .A4(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n831_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n710_), .A2(new_n386_), .A3(new_n723_), .A4(new_n274_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT118), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n639_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n843_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n343_), .A3(new_n614_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1340gat));
  NOR2_X1   g647(.A1(new_n574_), .A2(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n846_), .B1(KEYINPUT60), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n574_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G120gat), .B1(new_n852_), .B2(new_n844_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(KEYINPUT60), .B2(new_n850_), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n844_), .A2(new_n855_), .A3(new_n634_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G127gat), .B1(new_n846_), .B2(new_n647_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n858_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n856_), .B1(new_n859_), .B2(new_n860_), .ZN(G1342gat));
  OAI21_X1  g660(.A(G134gat), .B1(new_n844_), .B2(new_n646_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n846_), .A2(new_n528_), .A3(new_n536_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1343gat));
  NAND2_X1  g663(.A1(new_n840_), .A2(new_n448_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n865_), .A2(new_n651_), .A3(new_n274_), .A4(new_n660_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n614_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n851_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT120), .B(G148gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1345gat));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n647_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  NAND3_X1  g673(.A1(new_n866_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n866_), .A2(new_n692_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n530_), .ZN(G1347gat));
  OAI21_X1  g676(.A(new_n829_), .B1(new_n828_), .B2(new_n536_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n819_), .A2(new_n824_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(KEYINPUT57), .A3(new_n699_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n880_), .A3(new_n812_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n838_), .B1(new_n881_), .B2(new_n634_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n710_), .A2(new_n386_), .A3(new_n448_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n614_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n882_), .A2(new_n451_), .A3(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT121), .B1(new_n885_), .B2(new_n298_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n884_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n840_), .A2(new_n274_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(G169gat), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n886_), .A2(KEYINPUT62), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT121), .B(new_n892_), .C1(new_n885_), .C2(new_n298_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n885_), .A2(new_n311_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT122), .B1(new_n891_), .B2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n886_), .A2(new_n890_), .A3(KEYINPUT62), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n894_), .A4(new_n893_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1348gat));
  NOR2_X1   g699(.A1(new_n882_), .A2(new_n451_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n901_), .A2(new_n883_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n851_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT123), .B(G176gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1349gat));
  AND3_X1   g704(.A1(new_n901_), .A2(new_n647_), .A3(new_n883_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n396_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n906_), .B2(G183gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT124), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n908_), .B(new_n911_), .C1(G183gat), .C2(new_n906_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1350gat));
  NAND4_X1  g712(.A1(new_n902_), .A2(new_n393_), .A3(new_n395_), .A4(new_n536_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n902_), .A2(new_n692_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n288_), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n660_), .A2(new_n449_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n865_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(G197gat), .A3(new_n614_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n919_), .A2(KEYINPUT125), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(KEYINPUT125), .ZN(new_n921_));
  AOI21_X1  g720(.A(G197gat), .B1(new_n918_), .B2(new_n614_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(G1352gat));
  NAND2_X1  g722(.A1(new_n918_), .A2(new_n851_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n250_), .A2(KEYINPUT126), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1353gat));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n634_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n918_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n927_), .B1(new_n918_), .B2(new_n928_), .ZN(new_n931_));
  OAI22_X1  g730(.A1(new_n930_), .A2(new_n931_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n931_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n934_), .A3(new_n929_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n935_), .ZN(G1354gat));
  OR2_X1    g735(.A1(new_n865_), .A2(new_n917_), .ZN(new_n937_));
  OR3_X1    g736(.A1(new_n937_), .A2(G218gat), .A3(new_n699_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G218gat), .B1(new_n937_), .B2(new_n646_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1355gat));
endmodule


