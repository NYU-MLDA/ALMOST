//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_;
  XNOR2_X1  g000(.A(KEYINPUT10), .B(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G85gat), .B(G92gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(KEYINPUT9), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(KEYINPUT65), .A3(new_n212_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n208_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n207_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT8), .ZN(new_n225_));
  INV_X1    g024(.A(new_n209_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n206_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT6), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT6), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(KEYINPUT66), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(KEYINPUT6), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n206_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n226_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n228_), .B1(new_n240_), .B2(KEYINPUT67), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n225_), .B1(new_n238_), .B2(new_n226_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n217_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G36gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G29gat), .ZN(new_n247_));
  INV_X1    g046(.A(G29gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G36gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G50gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G43gat), .ZN(new_n252_));
  INV_X1    g051(.A(G43gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G50gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n245_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n215_), .A2(new_n216_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n208_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n237_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n209_), .B1(new_n263_), .B2(new_n234_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n264_), .A2(KEYINPUT67), .A3(new_n225_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n227_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n258_), .B(KEYINPUT15), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT34), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT35), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n259_), .A2(new_n269_), .A3(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n272_), .A2(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT72), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT36), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n276_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n259_), .A2(new_n269_), .A3(new_n284_), .A4(new_n274_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n277_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n281_), .B(new_n282_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n277_), .B2(new_n285_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n290_), .B1(KEYINPUT81), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(KEYINPUT81), .B2(new_n291_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT80), .B(G190gat), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n293_), .B(new_n294_), .C1(new_n291_), .C2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  INV_X1    g097(.A(G183gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT23), .B1(new_n299_), .B2(new_n290_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G183gat), .A3(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT82), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(KEYINPUT82), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n296_), .A2(new_n304_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(KEYINPUT83), .A3(new_n302_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n311_), .B(KEYINPUT23), .C1(new_n299_), .C2(new_n290_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n310_), .B(new_n312_), .C1(G183gat), .C2(new_n295_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G169gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(new_n253_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n317_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G127gat), .B(G134gat), .Z(new_n321_));
  XOR2_X1   g120(.A(G113gat), .B(G120gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n320_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G227gat), .A2(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(G15gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT30), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT31), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n324_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT92), .Z(new_n332_));
  INV_X1    g131(.A(G141gat), .ZN(new_n333_));
  INV_X1    g132(.A(G148gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(KEYINPUT84), .B2(KEYINPUT3), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT85), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT2), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(KEYINPUT85), .A3(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n336_), .A2(new_n339_), .A3(new_n341_), .A4(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n349_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n321_), .B(new_n322_), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n354_), .A2(new_n355_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n344_), .A2(new_n347_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(new_n323_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n360_), .B(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT91), .B1(new_n364_), .B2(KEYINPUT4), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n360_), .A2(new_n363_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n354_), .A2(new_n355_), .A3(new_n361_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT4), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT91), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n332_), .B(new_n359_), .C1(new_n365_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n332_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT93), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT0), .B(G57gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n382_), .B(KEYINPUT87), .Z(new_n383_));
  XNOR2_X1  g182(.A(G197gat), .B(G204gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT21), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT86), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n391_), .A3(new_n388_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n386_), .A2(new_n388_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n384_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(KEYINPUT21), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(G228gat), .A3(G233gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n401_), .A3(new_n398_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n383_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(new_n383_), .A3(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n407_));
  XOR2_X1   g206(.A(G22gat), .B(G50gat), .Z(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT28), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n403_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n404_), .A2(new_n411_), .A3(new_n405_), .A4(new_n410_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n379_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n381_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n397_), .A2(new_n317_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT26), .B(G190gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n294_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n306_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(KEYINPUT89), .A3(new_n306_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n310_), .A2(new_n312_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n298_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n303_), .B1(G183gat), .B2(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n315_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(KEYINPUT20), .B(new_n418_), .C1(new_n430_), .C2(new_n397_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT19), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n436_));
  INV_X1    g235(.A(new_n397_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n317_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n430_), .A2(new_n397_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n433_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT18), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n444_), .B(new_n445_), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n446_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n435_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n446_), .B(KEYINPUT97), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n426_), .A2(new_n298_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n424_), .B2(new_n423_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n429_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT95), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT95), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n427_), .A2(new_n459_), .A3(new_n429_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n460_), .A3(new_n437_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT96), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT20), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n418_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n461_), .B2(KEYINPUT20), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n433_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n439_), .A2(new_n434_), .A3(new_n440_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n454_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n453_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  AOI211_X1 g269(.A(KEYINPUT98), .B(new_n454_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n417_), .B(new_n452_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n415_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n373_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n364_), .A2(KEYINPUT91), .A3(KEYINPUT4), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n368_), .A2(new_n369_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n476_), .A2(new_n477_), .B1(new_n358_), .B2(new_n357_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n478_), .B2(new_n332_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT94), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(KEYINPUT33), .A4(new_n379_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n372_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n379_), .B1(new_n364_), .B2(new_n332_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n450_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n371_), .A2(KEYINPUT33), .A3(new_n373_), .A4(new_n379_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT94), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n380_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n481_), .A2(new_n484_), .A3(new_n486_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n466_), .A2(new_n467_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n446_), .A2(KEYINPUT32), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n442_), .A2(new_n491_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n493_), .B(new_n494_), .C1(new_n416_), .C2(new_n381_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n474_), .B1(new_n489_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n330_), .B1(new_n473_), .B2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n381_), .A2(new_n416_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(new_n330_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n470_), .A2(new_n471_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n415_), .A4(new_n452_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n289_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT12), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT68), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n509_));
  INV_X1    g308(.A(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n506_), .A2(KEYINPUT11), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n505_), .B(new_n508_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G57gat), .B(G64gat), .Z(new_n515_));
  INV_X1    g314(.A(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n505_), .B1(new_n518_), .B2(new_n508_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n504_), .B1(new_n245_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(G230gat), .ZN(new_n522_));
  INV_X1    g321(.A(G233gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n245_), .B2(new_n520_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n267_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT67), .B1(new_n264_), .B2(new_n225_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(new_n244_), .A3(new_n227_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT69), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n262_), .A4(new_n520_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n262_), .B(new_n520_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT69), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n520_), .B1(new_n531_), .B2(new_n262_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n524_), .B(new_n533_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G120gat), .B(G148gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n529_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n529_), .B2(new_n537_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT71), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT71), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G1gat), .A2(G8gat), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(KEYINPUT74), .A3(KEYINPUT14), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n326_), .A2(G22gat), .ZN(new_n554_));
  INV_X1    g353(.A(G22gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G15gat), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n553_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(G1gat), .A2(G8gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(G1gat), .A2(G8gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT75), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(G1gat), .ZN(new_n561_));
  INV_X1    g360(.A(G8gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n552_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT74), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n558_), .B2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n557_), .A2(new_n560_), .A3(new_n565_), .A4(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n553_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n560_), .A2(new_n565_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n518_), .A2(new_n508_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n578_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n576_), .A2(new_n577_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n520_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(new_n576_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n583_), .B(KEYINPUT17), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n576_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT76), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT76), .ZN(new_n594_));
  INV_X1    g393(.A(new_n257_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n247_), .A2(new_n249_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n593_), .A2(new_n597_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT77), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n569_), .A2(new_n573_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT76), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT76), .B1(new_n256_), .B2(new_n257_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n600_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n597_), .A2(new_n569_), .A3(new_n573_), .A4(new_n593_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT77), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n599_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT78), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n601_), .A2(new_n604_), .A3(new_n600_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n606_), .A2(KEYINPUT77), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(KEYINPUT78), .A3(new_n599_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G169gat), .B(G197gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(KEYINPUT79), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n268_), .A2(new_n574_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n615_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n611_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n617_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n621_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n551_), .A2(new_n592_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n503_), .A2(new_n631_), .A3(KEYINPUT100), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT100), .B1(new_n503_), .B2(new_n631_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n498_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT101), .Z(new_n637_));
  AOI21_X1  g436(.A(new_n630_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n551_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n289_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n642_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n592_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n638_), .A2(new_n639_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n561_), .A3(new_n499_), .A4(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT38), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n637_), .A2(new_n652_), .ZN(G1324gat));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n501_), .A2(new_n452_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n562_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n503_), .A2(new_n631_), .A3(new_n655_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n562_), .B1(KEYINPUT102), .B2(KEYINPUT39), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n658_), .A2(new_n657_), .A3(new_n659_), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n654_), .A2(new_n656_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g462(.A1(new_n503_), .A2(new_n631_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n330_), .B1(new_n666_), .B2(new_n632_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n326_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n330_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT41), .B1(new_n671_), .B2(G15gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n326_), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n669_), .A2(new_n672_), .B1(new_n654_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT103), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  OAI221_X1 g475(.A(new_n676_), .B1(new_n654_), .B2(new_n673_), .C1(new_n669_), .C2(new_n672_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n635_), .A2(new_n415_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n555_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(new_n681_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n474_), .A2(new_n555_), .ZN(new_n684_));
  OAI22_X1  g483(.A1(new_n682_), .A2(new_n683_), .B1(new_n654_), .B2(new_n684_), .ZN(G1327gat));
  NAND4_X1  g484(.A1(new_n638_), .A2(new_n289_), .A3(new_n592_), .A4(new_n639_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(G29gat), .A3(new_n498_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n592_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n551_), .A2(new_n688_), .A3(new_n630_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n497_), .A2(new_n502_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n645_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n644_), .C1(new_n497_), .C2(new_n502_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n689_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n499_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n687_), .B1(new_n698_), .B2(G29gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT105), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n696_), .A2(new_n655_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n655_), .A2(KEYINPUT106), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n655_), .A2(KEYINPUT106), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n686_), .A2(G36gat), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n702_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n702_), .B2(new_n709_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1329gat));
  NOR2_X1   g512(.A1(new_n330_), .A2(new_n253_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n696_), .A2(new_n697_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT109), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n696_), .A2(new_n717_), .A3(new_n697_), .A4(new_n714_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n253_), .B1(new_n686_), .B2(new_n330_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n716_), .A2(new_n722_), .A3(new_n718_), .A4(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  NAND4_X1  g523(.A1(new_n696_), .A2(G50gat), .A3(new_n474_), .A4(new_n697_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n251_), .B1(new_n686_), .B2(new_n415_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n629_), .A2(new_n592_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n503_), .A2(new_n551_), .A3(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n498_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n629_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(new_n551_), .A3(new_n646_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n499_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1332gat));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n705_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n733_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n729_), .A2(new_n705_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G64gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT48), .B(new_n737_), .C1(new_n729_), .C2(new_n705_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT111), .Z(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n729_), .B2(new_n670_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT49), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n733_), .A2(new_n747_), .A3(new_n670_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(new_n752_), .A3(new_n474_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n729_), .A2(new_n474_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G78gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT50), .B(new_n752_), .C1(new_n729_), .C2(new_n474_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT112), .Z(G1335gat));
  NOR3_X1   g558(.A1(new_n639_), .A2(new_n688_), .A3(new_n629_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n498_), .ZN(new_n762_));
  AND4_X1   g561(.A1(new_n289_), .A2(new_n732_), .A3(new_n592_), .A4(new_n551_), .ZN(new_n763_));
  INV_X1    g562(.A(G85gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n499_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1336gat));
  AOI21_X1  g565(.A(G92gat), .B1(new_n763_), .B2(new_n655_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT113), .Z(new_n768_));
  NOR3_X1   g567(.A1(new_n761_), .A2(new_n211_), .A3(new_n706_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1337gat));
  NAND3_X1  g569(.A1(new_n763_), .A2(new_n670_), .A3(new_n203_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n763_), .A2(new_n773_), .A3(new_n670_), .A4(new_n203_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n670_), .B(new_n760_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G99gat), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n776_), .A3(G99gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT51), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n775_), .B(new_n782_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1338gat));
  OAI211_X1 g583(.A(new_n474_), .B(new_n760_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(G106gat), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT52), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(G106gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n763_), .A2(new_n474_), .A3(new_n204_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n548_), .A2(new_n644_), .A3(new_n728_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT54), .ZN(new_n798_));
  INV_X1    g597(.A(new_n620_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT78), .B1(new_n615_), .B2(new_n599_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n609_), .B(new_n598_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n612_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n623_), .A2(new_n612_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n800_), .A2(new_n801_), .A3(new_n611_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n624_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n620_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n546_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n529_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT56), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n528_), .B1(new_n536_), .B2(KEYINPUT12), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n534_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n528_), .B(new_n534_), .C1(new_n536_), .C2(KEYINPUT12), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n524_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n521_), .A2(new_n525_), .A3(KEYINPUT55), .A4(new_n528_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n542_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n812_), .B1(new_n815_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n542_), .A3(new_n814_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n810_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT57), .B1(new_n827_), .B2(new_n289_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  INV_X1    g628(.A(new_n289_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n826_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n814_), .B1(new_n823_), .B2(new_n542_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n812_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n829_), .B(new_n830_), .C1(new_n833_), .C2(new_n810_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n823_), .A2(new_n835_), .A3(new_n542_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n824_), .A2(KEYINPUT56), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n610_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n620_), .B1(new_n838_), .B2(new_n803_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n799_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT118), .B1(new_n841_), .B2(new_n811_), .ZN(new_n842_));
  AND4_X1   g641(.A1(KEYINPUT118), .A2(new_n805_), .A3(new_n808_), .A4(new_n811_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n836_), .B(new_n837_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n644_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n809_), .B2(new_n544_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n841_), .A2(KEYINPUT118), .A3(new_n811_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT58), .A3(new_n836_), .A4(new_n837_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n828_), .A2(new_n834_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n592_), .B1(new_n852_), .B2(KEYINPUT119), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n828_), .A2(new_n834_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n846_), .A2(new_n851_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(KEYINPUT119), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n798_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n824_), .A2(new_n815_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(new_n629_), .A3(new_n811_), .A4(new_n826_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n810_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n829_), .B1(new_n863_), .B2(new_n830_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n827_), .A2(KEYINPUT57), .A3(new_n289_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n855_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n852_), .A2(KEYINPUT119), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n592_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(KEYINPUT120), .A3(new_n798_), .ZN(new_n871_));
  NOR4_X1   g670(.A1(new_n655_), .A2(new_n498_), .A3(new_n474_), .A4(new_n330_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n859_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n629_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n798_), .B1(new_n852_), .B2(new_n688_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n872_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n859_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n630_), .B(new_n879_), .C1(new_n880_), .C2(KEYINPUT59), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n875_), .B1(new_n881_), .B2(new_n874_), .ZN(G1340gat));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n884_));
  AOI21_X1  g683(.A(G120gat), .B1(new_n551_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n884_), .B2(G120gat), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n883_), .B1(new_n873_), .B2(new_n886_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n873_), .A2(new_n883_), .A3(new_n886_), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n639_), .B(new_n879_), .C1(new_n880_), .C2(KEYINPUT59), .ZN(new_n889_));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI22_X1  g689(.A1(new_n887_), .A2(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1341gat));
  NAND2_X1  g690(.A1(new_n688_), .A2(G127gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT122), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n879_), .B(new_n894_), .C1(new_n880_), .C2(KEYINPUT59), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n859_), .A2(new_n871_), .A3(new_n688_), .A4(new_n872_), .ZN(new_n896_));
  INV_X1    g695(.A(G127gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT123), .B1(new_n895_), .B2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n878_), .B(new_n893_), .C1(new_n873_), .C2(new_n877_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n898_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(G1342gat));
  INV_X1    g703(.A(G134gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n873_), .A2(new_n905_), .A3(new_n289_), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n644_), .B(new_n879_), .C1(new_n880_), .C2(KEYINPUT59), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n905_), .ZN(G1343gat));
  NAND2_X1  g707(.A1(new_n859_), .A2(new_n871_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n670_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n705_), .A2(new_n498_), .A3(new_n415_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(new_n333_), .A3(new_n629_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n911_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G141gat), .B1(new_n914_), .B2(new_n630_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1344gat));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n334_), .A3(new_n551_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G148gat), .B1(new_n914_), .B2(new_n639_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1345gat));
  XNOR2_X1  g718(.A(KEYINPUT61), .B(G155gat), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n912_), .A2(new_n688_), .A3(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n914_), .B2(new_n592_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1346gat));
  INV_X1    g723(.A(G162gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n644_), .A2(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT124), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n910_), .A2(new_n289_), .A3(new_n911_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n912_), .A2(new_n927_), .B1(new_n928_), .B2(new_n925_), .ZN(G1347gat));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n876_), .A2(new_n415_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n705_), .A2(new_n500_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n630_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT22), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n930_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(G169gat), .ZN(new_n937_));
  INV_X1    g736(.A(G169gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n934_), .B2(new_n930_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(new_n936_), .B2(new_n939_), .ZN(G1348gat));
  INV_X1    g739(.A(new_n933_), .ZN(new_n941_));
  AOI21_X1  g740(.A(G176gat), .B1(new_n941_), .B2(new_n551_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n909_), .A2(new_n474_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n932_), .A2(G176gat), .A3(new_n551_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n942_), .B1(new_n943_), .B2(new_n945_), .ZN(G1349gat));
  NAND3_X1  g745(.A1(new_n943_), .A2(new_n688_), .A3(new_n932_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n932_), .A2(new_n688_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n294_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n947_), .A2(new_n299_), .B1(new_n931_), .B2(new_n949_), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n933_), .B2(new_n644_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n289_), .A2(new_n419_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n933_), .B2(new_n952_), .ZN(G1351gat));
  AND2_X1   g752(.A1(new_n705_), .A2(new_n417_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n859_), .A2(new_n871_), .A3(new_n330_), .A4(new_n954_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n955_), .A2(new_n630_), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n956_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g756(.A1(new_n955_), .A2(new_n639_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n958_), .B(new_n959_), .ZN(G1353gat));
  NOR2_X1   g759(.A1(new_n955_), .A2(new_n592_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n961_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(KEYINPUT63), .B(G211gat), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n955_), .A2(new_n592_), .A3(new_n963_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n962_), .A2(new_n964_), .ZN(G1354gat));
  INV_X1    g764(.A(G218gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n966_), .B1(new_n955_), .B2(new_n830_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n857_), .A2(new_n858_), .ZN(new_n968_));
  AOI21_X1  g767(.A(KEYINPUT120), .B1(new_n870_), .B2(new_n798_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n644_), .A2(new_n966_), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n971_), .B(KEYINPUT126), .ZN(new_n972_));
  NAND4_X1  g771(.A1(new_n970_), .A2(new_n330_), .A3(new_n954_), .A4(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n967_), .A2(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(new_n975_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n967_), .A2(new_n973_), .A3(KEYINPUT127), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1355gat));
endmodule


