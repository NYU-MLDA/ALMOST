//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  OR3_X1    g011(.A1(new_n211_), .A2(KEYINPUT89), .A3(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT89), .B1(new_n211_), .B2(new_n212_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT87), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n219_), .A2(KEYINPUT87), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n217_), .B(new_n218_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n211_), .A2(new_n215_), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n219_), .B(KEYINPUT3), .Z(new_n224_));
  XOR2_X1   g023(.A(new_n218_), .B(KEYINPUT2), .Z(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n227_), .A2(new_n231_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(KEYINPUT4), .ZN(new_n238_));
  INV_X1    g037(.A(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(KEYINPUT96), .A3(KEYINPUT4), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n222_), .A2(new_n226_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n230_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n237_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT96), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n240_), .B1(new_n241_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT97), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n236_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n241_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n240_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n250_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n206_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT97), .ZN(new_n255_));
  INV_X1    g054(.A(new_n206_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n247_), .A2(new_n248_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .A4(new_n236_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT98), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n262_));
  OR3_X1    g061(.A1(new_n227_), .A2(KEYINPUT29), .A3(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G22gat), .B(G50gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G211gat), .B(G218gat), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(G197gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(G197gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT21), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n270_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT91), .B1(new_n270_), .B2(G197gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n269_), .B(new_n273_), .C1(new_n276_), .C2(KEYINPUT21), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n269_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n242_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G228gat), .ZN(new_n284_));
  INV_X1    g083(.A(G233gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n281_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G78gat), .B(G106gat), .Z(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT92), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n290_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n291_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT93), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n297_));
  AOI211_X1 g096(.A(new_n297_), .B(new_n291_), .C1(new_n287_), .C2(new_n290_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n268_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n268_), .A2(new_n292_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n291_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n253_), .A2(new_n258_), .A3(KEYINPUT98), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT23), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(G183gat), .B2(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT22), .B(G169gat), .Z(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(new_n312_), .C1(G176gat), .C2(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n312_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n318_), .B(new_n310_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n322_), .A2(new_n281_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT94), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT19), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n288_), .A2(new_n321_), .A3(new_n314_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT20), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n326_), .B1(new_n329_), .B2(new_n323_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n331_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n308_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n329_), .A2(new_n326_), .A3(new_n323_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n324_), .A2(new_n330_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(new_n326_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT27), .B(new_n338_), .C1(new_n344_), .C2(new_n336_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n261_), .A2(new_n306_), .A3(new_n307_), .A4(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n339_), .A2(new_n340_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n250_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n234_), .A2(new_n239_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n206_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n349_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT33), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n353_), .B1(new_n258_), .B2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n249_), .A2(new_n252_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(KEYINPUT33), .A3(new_n256_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n331_), .A2(new_n337_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n336_), .A2(KEYINPUT32), .ZN(new_n359_));
  MUX2_X1   g158(.A(new_n344_), .B(new_n358_), .S(new_n359_), .Z(new_n360_));
  AOI22_X1  g159(.A1(new_n355_), .A2(new_n357_), .B1(new_n259_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n348_), .B1(new_n361_), .B2(new_n306_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n322_), .B(KEYINPUT30), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(new_n230_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G99gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n365_), .B(new_n231_), .ZN(new_n368_));
  INV_X1    g167(.A(G99gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT86), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT83), .B(KEYINPUT84), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G71gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n375_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n371_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n367_), .A2(new_n370_), .A3(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n253_), .A2(KEYINPUT98), .A3(new_n258_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT98), .B1(new_n253_), .B2(new_n258_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n300_), .A2(new_n304_), .A3(new_n346_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(KEYINPUT100), .A3(new_n382_), .A4(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n261_), .A2(new_n307_), .A3(new_n387_), .A4(new_n382_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT100), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n362_), .A2(new_n383_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G106gat), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n369_), .A2(KEYINPUT10), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n369_), .A2(KEYINPUT10), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G99gat), .A2(G106gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G85gat), .A2(G92gat), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n402_), .A2(KEYINPUT9), .ZN(new_n403_));
  INV_X1    g202(.A(G92gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n203_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT9), .A3(new_n402_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n396_), .A2(new_n401_), .A3(new_n403_), .A4(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT7), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n369_), .A3(new_n393_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n409_), .A2(new_n399_), .A3(new_n400_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT8), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n405_), .A2(new_n402_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n407_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G57gat), .ZN(new_n417_));
  INV_X1    g216(.A(G64gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G57gat), .A2(G64gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT11), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G71gat), .B(G78gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT11), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n419_), .A2(new_n425_), .A3(new_n420_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n423_), .A3(KEYINPUT11), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n416_), .A2(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n429_), .B(new_n407_), .C1(new_n415_), .C2(new_n414_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G230gat), .A2(G233gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(KEYINPUT64), .Z(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G120gat), .B(G148gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT68), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT67), .Z(new_n441_));
  XOR2_X1   g240(.A(G176gat), .B(G204gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT5), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n441_), .B(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n431_), .A2(KEYINPUT12), .A3(new_n432_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n416_), .A2(new_n446_), .A3(new_n430_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n435_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT66), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451_));
  AOI211_X1 g250(.A(new_n451_), .B(new_n435_), .C1(new_n445_), .C2(new_n447_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n438_), .B(new_n444_), .C1(new_n450_), .C2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n436_), .B(KEYINPUT65), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n449_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n451_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n435_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT66), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n454_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n444_), .B(KEYINPUT69), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n453_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT13), .ZN(new_n464_));
  OAI211_X1 g263(.A(KEYINPUT70), .B(new_n453_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n464_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n469_), .A2(KEYINPUT71), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(KEYINPUT71), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G1gat), .A2(G8gat), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n474_), .A2(KEYINPUT77), .A3(KEYINPUT14), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT77), .B1(new_n474_), .B2(KEYINPUT14), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT78), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT78), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n479_), .B(new_n473_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G1gat), .B(G8gat), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n478_), .A2(new_n482_), .A3(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G29gat), .B(G36gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT15), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n492_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n485_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n482_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n489_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n489_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n495_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n494_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT82), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n494_), .A2(new_n501_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n509_), .B2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n472_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n392_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n490_), .A2(new_n416_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n416_), .A2(new_n498_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G232gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT34), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n515_), .B(new_n516_), .C1(KEYINPUT35), .C2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT35), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT72), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n519_), .B(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G190gat), .B(G218gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT74), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT75), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n532_), .B1(new_n533_), .B2(KEYINPUT37), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(KEYINPUT37), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT76), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n534_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n486_), .A2(G231gat), .A3(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n484_), .A2(new_n485_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n429_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n430_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G211gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT16), .B(G183gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT79), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n551_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n540_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n540_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT80), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT80), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n547_), .A2(new_n551_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n554_), .B2(new_n551_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n557_), .B(new_n560_), .C1(new_n562_), .C2(new_n540_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n539_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n514_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OR3_X1    g366(.A1(new_n567_), .A2(G1gat), .A3(new_n386_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n569_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n556_), .A2(new_n558_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n532_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n514_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G1gat), .B1(new_n575_), .B2(new_n386_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n571_), .A3(new_n576_), .ZN(G1324gat));
  INV_X1    g376(.A(G8gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n566_), .A2(new_n578_), .A3(new_n346_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n348_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n355_), .A2(new_n357_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n259_), .A2(new_n360_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n306_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n383_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n388_), .A2(new_n391_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n513_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n346_), .A4(new_n574_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT102), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n578_), .B1(new_n588_), .B2(KEYINPUT102), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n579_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(G1325gat));
  OR3_X1    g395(.A1(new_n567_), .A2(G15gat), .A3(new_n383_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G15gat), .B1(new_n575_), .B2(new_n383_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT41), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT41), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(G1326gat));
  INV_X1    g400(.A(new_n306_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G22gat), .B1(new_n575_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT42), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n602_), .A2(G22gat), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n604_), .B1(new_n567_), .B2(new_n605_), .ZN(G1327gat));
  INV_X1    g405(.A(new_n564_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n532_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n514_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(G29gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n386_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n513_), .B1(KEYINPUT104), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n586_), .B2(new_n539_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT43), .B(new_n538_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n564_), .B(new_n615_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n614_), .A2(KEYINPUT104), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n392_), .B2(new_n538_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n586_), .A2(new_n616_), .A3(new_n539_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n607_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n620_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n615_), .A3(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n386_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n613_), .B1(new_n627_), .B2(new_n611_), .ZN(G1328gat));
  NAND2_X1  g427(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n623_), .ZN(new_n630_));
  AND4_X1   g429(.A1(new_n564_), .A2(new_n630_), .A3(new_n615_), .A4(new_n625_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n625_), .B1(new_n624_), .B2(new_n615_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n346_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n635_));
  INV_X1    g434(.A(G36gat), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n514_), .A2(new_n636_), .A3(new_n346_), .A4(new_n608_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT45), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT45), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n629_), .B1(new_n634_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n347_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n629_), .B(new_n640_), .C1(new_n642_), .C2(new_n636_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n644_), .ZN(G1329gat));
  NOR3_X1   g444(.A1(new_n609_), .A2(G43gat), .A3(new_n383_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n383_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n648_));
  INV_X1    g447(.A(G43gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT47), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT47), .B(new_n647_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1330gat));
  INV_X1    g453(.A(G50gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n610_), .A2(new_n655_), .A3(new_n306_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n602_), .B1(new_n621_), .B2(new_n626_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(new_n655_), .ZN(G1331gat));
  NOR2_X1   g457(.A1(new_n472_), .A2(new_n512_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n586_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n564_), .A2(new_n573_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n662_), .A2(new_n417_), .A3(new_n386_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n565_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n612_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n663_), .B1(new_n417_), .B2(new_n666_), .ZN(G1332gat));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n418_), .A3(new_n346_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G64gat), .B1(new_n662_), .B2(new_n347_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n672_), .B2(new_n673_), .ZN(G1333gat));
  OR3_X1    g473(.A1(new_n664_), .A2(G71gat), .A3(new_n383_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n660_), .A2(new_n382_), .A3(new_n661_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT49), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G71gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G71gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT107), .ZN(G1334gat));
  OAI21_X1  g480(.A(G78gat), .B1(new_n662_), .B2(new_n602_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT50), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n602_), .A2(G78gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n664_), .B2(new_n684_), .ZN(G1335gat));
  NAND2_X1  g484(.A1(new_n660_), .A2(new_n608_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G85gat), .B1(new_n687_), .B2(new_n612_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n624_), .A2(new_n659_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n386_), .A2(new_n203_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(G1336gat));
  OAI21_X1  g490(.A(new_n404_), .B1(new_n686_), .B2(new_n347_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n692_), .A2(new_n693_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n347_), .A2(new_n404_), .ZN(new_n696_));
  AOI211_X1 g495(.A(new_n694_), .B(new_n695_), .C1(new_n689_), .C2(new_n696_), .ZN(G1337gat));
  OAI21_X1  g496(.A(new_n382_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n686_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n689_), .A2(new_n382_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G99gat), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1338gat));
  NAND3_X1  g502(.A1(new_n687_), .A2(new_n393_), .A3(new_n306_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n624_), .A2(new_n306_), .A3(new_n659_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G106gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G106gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT53), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT53), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1339gat));
  INV_X1    g512(.A(KEYINPUT116), .ZN(new_n714_));
  INV_X1    g513(.A(new_n572_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n512_), .A2(new_n453_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n460_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT55), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n445_), .A2(new_n435_), .A3(new_n447_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(KEYINPUT55), .B2(new_n457_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n719_), .B2(new_n722_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n717_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT56), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT56), .B(new_n717_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n716_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n491_), .A2(new_n495_), .A3(new_n493_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n492_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n504_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(KEYINPUT111), .A3(new_n504_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT112), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n498_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n495_), .B1(new_n738_), .B2(new_n493_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n734_), .B1(new_n739_), .B2(new_n505_), .ZN(new_n740_));
  AND4_X1   g539(.A1(KEYINPUT112), .A2(new_n740_), .A3(new_n736_), .A4(new_n730_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n507_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT113), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n507_), .C1(new_n737_), .C2(new_n741_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n743_), .A2(new_n745_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n532_), .B1(new_n729_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT57), .B(new_n532_), .C1(new_n729_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT55), .B1(new_n456_), .B2(new_n458_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n457_), .A2(KEYINPUT55), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n449_), .B2(new_n448_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n719_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n460_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n759_), .B2(KEYINPUT56), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n725_), .A2(KEYINPUT114), .A3(new_n726_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n728_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n743_), .A2(new_n745_), .B1(new_n459_), .B2(new_n444_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(KEYINPUT58), .A3(new_n763_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n539_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n751_), .B1(new_n752_), .B2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n538_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT115), .A3(new_n767_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n715_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773_));
  INV_X1    g572(.A(new_n512_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n559_), .A2(new_n563_), .A3(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n469_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n538_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n469_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT54), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n468_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n775_), .B1(new_n780_), .B2(new_n466_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT109), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n538_), .A4(new_n776_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n779_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n714_), .B1(new_n772_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n784_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n770_), .A2(KEYINPUT115), .A3(new_n767_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n770_), .B2(new_n767_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n751_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT116), .B(new_n787_), .C1(new_n790_), .C2(new_n715_), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n386_), .A2(new_n306_), .A3(new_n346_), .A4(new_n383_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n786_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n786_), .A2(new_n791_), .A3(KEYINPUT117), .A4(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n512_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(G113gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n749_), .A2(new_n750_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n607_), .B1(new_n802_), .B2(new_n768_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n804_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n787_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n792_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n774_), .A2(new_n800_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n793_), .A2(new_n811_), .A3(KEYINPUT59), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n793_), .B2(KEYINPUT59), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n809_), .B(new_n810_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n774_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(new_n815_), .B2(G113gat), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n801_), .A2(new_n814_), .A3(new_n816_), .ZN(G1340gat));
  INV_X1    g616(.A(new_n472_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n809_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G120gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n472_), .A2(KEYINPUT60), .ZN(new_n821_));
  MUX2_X1   g620(.A(new_n821_), .B(KEYINPUT60), .S(G120gat), .Z(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT121), .B1(new_n797_), .B2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n797_), .A2(KEYINPUT121), .A3(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n823_), .B2(new_n824_), .ZN(G1341gat));
  AOI21_X1  g624(.A(G127gat), .B1(new_n797_), .B2(new_n607_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n812_), .A2(new_n813_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n809_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n715_), .A2(G127gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n826_), .B1(new_n829_), .B2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n797_), .B2(new_n573_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n539_), .A2(G134gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n829_), .B2(new_n833_), .ZN(G1343gat));
  AND2_X1   g633(.A1(new_n786_), .A2(new_n791_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n612_), .A2(new_n306_), .A3(new_n347_), .A4(new_n383_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT122), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n512_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n472_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT123), .B(G148gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n838_), .A2(new_n564_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  AOI21_X1  g646(.A(G162gat), .B1(new_n839_), .B2(new_n573_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n539_), .A2(G162gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n839_), .B2(new_n849_), .ZN(G1347gat));
  NAND3_X1  g649(.A1(new_n386_), .A2(new_n346_), .A3(new_n382_), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n851_), .B(KEYINPUT124), .Z(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n306_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n807_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n512_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n313_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(G169gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n858_), .B2(new_n859_), .ZN(G1348gat));
  AOI21_X1  g660(.A(G176gat), .B1(new_n855_), .B2(new_n818_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n835_), .A2(new_n602_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n852_), .A2(G176gat), .A3(new_n818_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1349gat));
  NAND2_X1  g664(.A1(new_n807_), .A2(new_n854_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(new_n316_), .A3(new_n572_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n863_), .A2(new_n607_), .A3(new_n852_), .ZN(new_n870_));
  INV_X1    g669(.A(G183gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1350gat));
  OAI21_X1  g671(.A(G190gat), .B1(new_n866_), .B2(new_n538_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n573_), .A2(new_n317_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(KEYINPUT126), .Z(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n866_), .B2(new_n875_), .ZN(G1351gat));
  NOR4_X1   g675(.A1(new_n612_), .A2(new_n602_), .A3(new_n347_), .A4(new_n382_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n835_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n774_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT127), .B(G197gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1352gat));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n472_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(new_n270_), .ZN(G1353gat));
  AND2_X1   g682(.A1(new_n835_), .A2(new_n877_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n572_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n886_), .B(new_n887_), .Z(G1354gat));
  AOI21_X1  g687(.A(G218gat), .B1(new_n884_), .B2(new_n573_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n539_), .A2(G218gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n884_), .B2(new_n890_), .ZN(G1355gat));
endmodule


