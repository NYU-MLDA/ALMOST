//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT65), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(KEYINPUT65), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(new_n203_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT9), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n218_));
  OR2_X1    g017(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT64), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n223_), .A3(new_n220_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n213_), .B(new_n218_), .C1(new_n225_), .C2(G106gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n210_), .A2(new_n211_), .A3(new_n203_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n203_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT66), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n217_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT66), .B1(new_n213_), .B2(new_n230_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n229_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n227_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n228_), .B2(new_n229_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n241_), .B(new_n242_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n234_), .B1(new_n243_), .B2(new_n217_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n226_), .B1(new_n238_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT68), .B(new_n226_), .C1(new_n238_), .C2(new_n244_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G57gat), .B(G64gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(KEYINPUT11), .ZN(new_n251_));
  XOR2_X1   g050(.A(G71gat), .B(G78gat), .Z(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(new_n248_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n255_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n256_), .B(new_n258_), .C1(new_n259_), .C2(KEYINPUT12), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT69), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n247_), .A2(new_n248_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n257_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n256_), .A2(new_n258_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .A4(new_n261_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n263_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n256_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n262_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G120gat), .B(G148gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G176gat), .B(G204gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n273_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT13), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(KEYINPUT13), .A3(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G29gat), .B(G36gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G43gat), .B(G50gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT15), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n289_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G229gat), .A2(G233gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT76), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n296_), .B(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n301_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n300_), .A2(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G113gat), .B(G141gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(G169gat), .B(G197gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT77), .Z(new_n310_));
  OR2_X1    g109(.A1(new_n305_), .A2(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n286_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT22), .B(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT94), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G176gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT95), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n324_), .B(KEYINPUT79), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(new_n326_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n323_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n324_), .B(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT23), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT95), .B(new_n332_), .C1(new_n335_), .C2(new_n327_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n322_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT96), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT78), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT25), .B(G183gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n340_), .A2(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n325_), .A2(KEYINPUT81), .A3(new_n326_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n324_), .B2(KEYINPUT23), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n345_), .B(new_n347_), .C1(new_n328_), .C2(new_n326_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n339_), .B(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(KEYINPUT24), .A3(new_n316_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n344_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT93), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n344_), .A2(new_n348_), .A3(KEYINPUT93), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G197gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(G204gat), .ZN(new_n358_));
  INV_X1    g157(.A(G204gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(G197gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT21), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n358_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n363_), .B2(new_n358_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT89), .B(KEYINPUT21), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n361_), .B(new_n362_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n362_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT96), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n322_), .A2(new_n331_), .A3(new_n336_), .A4(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n338_), .A2(new_n356_), .A3(new_n371_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT19), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n348_), .A2(new_n332_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n321_), .A2(KEYINPUT80), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n321_), .B1(KEYINPUT80), .B2(KEYINPUT22), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n318_), .A2(new_n380_), .B1(G169gat), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n344_), .A2(new_n351_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n329_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n378_), .B1(new_n385_), .B2(new_n370_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n374_), .A2(new_n377_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n385_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n378_), .B1(new_n389_), .B2(new_n371_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n338_), .A2(new_n356_), .A3(new_n373_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n391_), .A2(KEYINPUT97), .A3(new_n370_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT97), .B1(new_n391_), .B2(new_n370_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n388_), .B1(new_n394_), .B2(new_n376_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT18), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  NOR2_X1   g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n399_), .ZN(new_n401_));
  AOI211_X1 g200(.A(new_n401_), .B(new_n388_), .C1(new_n394_), .C2(new_n376_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n315_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n386_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n371_), .A2(new_n337_), .A3(new_n352_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n376_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n394_), .B2(new_n376_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n401_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n395_), .A2(new_n399_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT27), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n403_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT98), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT83), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G141gat), .A3(G148gat), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G141gat), .ZN(new_n422_));
  INV_X1    g221(.A(G148gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n417_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT84), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n417_), .A2(new_n426_), .A3(new_n429_), .A4(new_n421_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT2), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n414_), .A2(new_n416_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT85), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n413_), .A2(new_n432_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n424_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n422_), .A2(new_n423_), .A3(KEYINPUT3), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n414_), .A2(new_n416_), .A3(new_n440_), .A4(new_n432_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n434_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n418_), .A2(new_n420_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n431_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(G127gat), .B(G134gat), .Z(new_n447_));
  XOR2_X1   g246(.A(G113gat), .B(G120gat), .Z(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n428_), .A2(new_n430_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n450_), .A2(new_n453_), .A3(KEYINPUT4), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(new_n455_), .A3(new_n449_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G225gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n412_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n450_), .A2(new_n453_), .A3(KEYINPUT4), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(KEYINPUT98), .A3(new_n458_), .A4(new_n456_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n450_), .A2(new_n453_), .A3(new_n457_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT99), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(G85gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT0), .B(G57gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n467_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n463_), .A2(new_n471_), .A3(new_n466_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT102), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT102), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n467_), .A2(new_n476_), .A3(new_n472_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n411_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n385_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n385_), .A2(new_n484_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G227gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(G15gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT30), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n481_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT82), .A3(new_n491_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n449_), .B(KEYINPUT31), .Z(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n481_), .B(new_n499_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n367_), .A2(new_n369_), .B1(G228gat), .B2(G233gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n431_), .B2(new_n445_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n504_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n451_), .A2(KEYINPUT87), .A3(new_n505_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT90), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n507_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT87), .B1(new_n451_), .B2(new_n505_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT90), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .A4(new_n504_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(G228gat), .B(G233gat), .C1(new_n371_), .C2(new_n506_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT28), .B1(new_n446_), .B2(KEYINPUT29), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n451_), .A2(new_n522_), .A3(new_n505_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G22gat), .B(G50gat), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n521_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n525_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n520_), .A2(new_n523_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT86), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n531_), .B2(new_n524_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n518_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n515_), .A2(KEYINPUT91), .A3(new_n516_), .A4(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n519_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n515_), .A2(new_n516_), .A3(new_n534_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n503_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n534_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n542_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n543_), .A2(KEYINPUT92), .A3(new_n539_), .A4(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n533_), .B1(new_n519_), .B2(new_n537_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n502_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  AOI211_X1 g347(.A(new_n501_), .B(new_n546_), .C1(new_n541_), .C2(new_n544_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n480_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n474_), .A2(KEYINPUT100), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT33), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n463_), .A2(new_n553_), .A3(new_n471_), .A4(new_n466_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT101), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n400_), .A2(new_n402_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n474_), .A2(new_n552_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n461_), .A2(new_n457_), .A3(new_n456_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n450_), .A2(new_n453_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n471_), .B1(new_n561_), .B2(new_n458_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT101), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n551_), .A2(new_n564_), .A3(new_n552_), .A4(new_n554_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n556_), .A2(new_n557_), .A3(new_n563_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n395_), .B1(new_n567_), .B2(new_n401_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n407_), .A2(KEYINPUT32), .A3(new_n399_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n475_), .A2(new_n568_), .A3(new_n569_), .A4(new_n477_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n545_), .A2(new_n501_), .A3(new_n547_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n550_), .A2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n314_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n247_), .A2(new_n289_), .A3(new_n248_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n578_), .A2(new_n579_), .B1(new_n245_), .B2(new_n290_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT70), .B1(new_n264_), .B2(new_n298_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT35), .Z(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n580_), .A2(new_n581_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(KEYINPUT35), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n577_), .B(new_n585_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(KEYINPUT73), .A3(new_n584_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT36), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n588_), .A2(KEYINPUT74), .A3(new_n589_), .A4(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n592_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT71), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT72), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n602_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n576_), .B(new_n594_), .C1(new_n597_), .C2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(KEYINPUT37), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n255_), .B(new_n296_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611_));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n610_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(KEYINPUT17), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n610_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n607_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n575_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT103), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(KEYINPUT103), .ZN(new_n624_));
  AND4_X1   g423(.A1(new_n202_), .A2(new_n623_), .A3(new_n479_), .A4(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT38), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT38), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n594_), .B1(new_n597_), .B2(new_n603_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n550_), .B2(new_n573_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT104), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT104), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR4_X1   g431(.A1(new_n632_), .A2(new_n620_), .A3(new_n313_), .A4(new_n286_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n202_), .B1(new_n633_), .B2(new_n479_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n626_), .A2(new_n627_), .A3(new_n634_), .ZN(G1324gat));
  NAND4_X1  g434(.A1(new_n623_), .A2(new_n292_), .A3(new_n411_), .A4(new_n624_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n286_), .A2(new_n620_), .A3(new_n313_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n411_), .B(new_n637_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(new_n639_), .A3(G8gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n638_), .B2(G8gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g442(.A1(new_n633_), .A2(new_n502_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n645_));
  AND3_X1   g444(.A1(new_n644_), .A2(G15gat), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n644_), .B2(G15gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n502_), .A2(new_n488_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n646_), .A2(new_n647_), .B1(new_n622_), .B2(new_n648_), .ZN(G1326gat));
  NAND2_X1  g448(.A1(new_n545_), .A2(new_n547_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OR3_X1    g450(.A1(new_n622_), .A2(G22gat), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n633_), .A2(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G22gat), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(new_n620_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n286_), .A2(new_n658_), .A3(new_n313_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n574_), .A2(new_n660_), .A3(new_n607_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n574_), .B2(new_n607_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n659_), .B(KEYINPUT44), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n478_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n628_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n658_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n575_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n478_), .A2(G29gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT106), .Z(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n671_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(new_n411_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT108), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(KEYINPUT108), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n671_), .A2(G36gat), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT45), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n665_), .A2(new_n411_), .A3(new_n666_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT107), .B1(new_n682_), .B2(G36gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n681_), .B(KEYINPUT46), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NOR2_X1   g488(.A1(new_n501_), .A2(new_n483_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n665_), .A2(new_n666_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n665_), .A2(KEYINPUT109), .A3(new_n666_), .A4(new_n690_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n483_), .B1(new_n671_), .B2(new_n501_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n693_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1330gat));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n667_), .A2(new_n699_), .A3(new_n651_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n575_), .A2(new_n650_), .A3(new_n670_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n699_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n286_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n312_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(new_n574_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n621_), .ZN(new_n706_));
  INV_X1    g505(.A(G57gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n479_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n704_), .A2(new_n658_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n632_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n479_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n712_), .B2(new_n707_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n714_), .A3(new_n678_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n709_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n678_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(G64gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(G64gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT111), .Z(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n710_), .B2(new_n502_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT49), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n706_), .A2(new_n723_), .A3(new_n502_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n710_), .B2(new_n650_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT50), .Z(new_n730_));
  NAND2_X1  g529(.A1(new_n650_), .A2(new_n728_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n706_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1335gat));
  OR2_X1    g533(.A1(new_n661_), .A2(new_n662_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n736_));
  OR3_X1    g535(.A1(new_n661_), .A2(new_n662_), .A3(KEYINPUT113), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n736_), .A2(new_n620_), .A3(new_n704_), .A4(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n478_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n705_), .A2(new_n670_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n214_), .A3(new_n479_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT114), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1336gat));
  OAI21_X1  g545(.A(G92gat), .B1(new_n738_), .B2(new_n679_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n215_), .A3(new_n411_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(KEYINPUT115), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n738_), .B2(new_n501_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n225_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n740_), .A2(new_n755_), .A3(new_n502_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1338gat));
  INV_X1    g560(.A(G106gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n740_), .A2(new_n762_), .A3(new_n650_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  NOR4_X1   g563(.A1(new_n703_), .A2(new_n651_), .A3(new_n658_), .A4(new_n312_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n735_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(G106gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT52), .B(new_n762_), .C1(new_n735_), .C2(new_n765_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g569(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n313_), .A2(new_n658_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n703_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n772_), .B1(new_n775_), .B2(new_n607_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n607_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(new_n703_), .A3(new_n774_), .A4(new_n771_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n263_), .A2(new_n780_), .A3(new_n270_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT118), .A4(new_n262_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n262_), .A2(KEYINPUT118), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n260_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n261_), .A2(new_n780_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n781_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n278_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT120), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n278_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n787_), .A2(new_n793_), .A3(KEYINPUT56), .A4(new_n278_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n297_), .A2(new_n299_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n302_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n797_), .B2(new_n796_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n308_), .B1(new_n303_), .B2(new_n302_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n310_), .A2(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n281_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n795_), .A2(KEYINPUT58), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n795_), .A2(new_n803_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n795_), .A2(KEYINPUT122), .A3(KEYINPUT58), .A4(new_n803_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n806_), .A2(new_n809_), .A3(new_n607_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n281_), .A2(new_n312_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n792_), .B2(new_n788_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n282_), .A2(new_n802_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n669_), .B(KEYINPUT57), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n813_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n628_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n811_), .A2(new_n815_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n779_), .B1(new_n620_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n675_), .A2(new_n549_), .A3(new_n479_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n815_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n811_), .A2(new_n818_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(KEYINPUT124), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT124), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n811_), .A2(new_n826_), .A3(new_n818_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n658_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n779_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT59), .B1(new_n821_), .B2(KEYINPUT123), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(KEYINPUT123), .B2(new_n821_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n312_), .B(new_n822_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G113gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n820_), .A2(new_n821_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n312_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(G1340gat));
  OAI211_X1 g636(.A(new_n286_), .B(new_n822_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n703_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n834_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(G1341gat));
  OAI211_X1 g642(.A(new_n658_), .B(new_n822_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G127gat), .ZN(new_n845_));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n834_), .A2(new_n846_), .A3(new_n658_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1342gat));
  OAI211_X1 g647(.A(new_n607_), .B(new_n822_), .C1(new_n829_), .C2(new_n831_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G134gat), .ZN(new_n850_));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n834_), .A2(new_n851_), .A3(new_n628_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1343gat));
  INV_X1    g652(.A(new_n548_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n819_), .A2(new_n620_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n776_), .A2(new_n778_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n679_), .A2(new_n479_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n858_), .A2(new_n313_), .A3(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n422_), .ZN(G1344gat));
  NOR3_X1   g660(.A1(new_n858_), .A2(new_n703_), .A3(new_n859_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n423_), .ZN(G1345gat));
  NAND4_X1  g662(.A1(new_n857_), .A2(new_n479_), .A3(new_n658_), .A4(new_n679_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  OR4_X1    g665(.A1(G162gat), .A2(new_n858_), .A3(new_n669_), .A4(new_n859_), .ZN(new_n867_));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n858_), .A2(new_n777_), .A3(new_n859_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n679_), .A2(new_n479_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n502_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n650_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n312_), .B(new_n873_), .C1(new_n828_), .C2(new_n779_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G169gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n825_), .A2(new_n827_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n856_), .B1(new_n879_), .B2(new_n658_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n880_), .A2(new_n320_), .A3(new_n312_), .A4(new_n873_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(new_n878_), .A3(new_n881_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n286_), .A3(new_n873_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n820_), .A2(new_n650_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n872_), .A2(new_n321_), .A3(new_n703_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n321_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n620_), .A2(new_n342_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n880_), .A2(new_n887_), .A3(new_n873_), .A4(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n872_), .A2(new_n620_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n884_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(G183gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n873_), .B(new_n888_), .C1(new_n828_), .C2(new_n779_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT125), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n889_), .A2(new_n893_), .A3(new_n895_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n880_), .A2(new_n607_), .A3(new_n873_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G190gat), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n880_), .A2(new_n628_), .A3(new_n343_), .A4(new_n873_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1351gat));
  AND2_X1   g699(.A1(new_n857_), .A2(new_n871_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n312_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n286_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT126), .B(G204gat), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n904_), .B(new_n906_), .ZN(G1353gat));
  NAND2_X1  g706(.A1(new_n855_), .A2(new_n856_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n620_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n908_), .A2(new_n548_), .A3(new_n871_), .A4(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT127), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n857_), .A2(new_n913_), .A3(new_n871_), .A4(new_n909_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n912_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n912_), .B1(new_n911_), .B2(new_n914_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1354gat));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n901_), .A2(new_n918_), .A3(new_n628_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n901_), .A2(new_n607_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n918_), .ZN(G1355gat));
endmodule


