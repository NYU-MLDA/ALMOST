//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G92gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(new_n203_), .A3(G85gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT9), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n204_), .A2(new_n207_), .A3(new_n210_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT66), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT66), .B1(new_n212_), .B2(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  INV_X1    g019(.A(G99gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n206_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n218_), .A2(new_n219_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(new_n209_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n208_), .A2(KEYINPUT65), .A3(new_n209_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT8), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n231_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n212_), .A2(new_n214_), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n233_), .B(new_n234_), .C1(new_n235_), .C2(new_n224_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n217_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G64gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n240_));
  XOR2_X1   g039(.A(G71gat), .B(G78gat), .Z(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n237_), .A2(new_n238_), .A3(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(KEYINPUT67), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n215_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT66), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n222_), .A2(new_n223_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n234_), .B1(new_n252_), .B2(new_n233_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n235_), .A2(new_n224_), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n254_), .A2(KEYINPUT8), .A3(new_n231_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n216_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n247_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n247_), .A2(new_n256_), .ZN(new_n258_));
  AOI211_X1 g057(.A(new_n246_), .B(new_n257_), .C1(new_n238_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n247_), .A2(new_n256_), .ZN(new_n262_));
  OAI211_X1 g061(.A(G230gat), .B(G233gat), .C1(new_n262_), .C2(new_n257_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G120gat), .B(G148gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT13), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(KEYINPUT13), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT89), .ZN(new_n279_));
  OR2_X1    g078(.A1(G197gat), .A2(G204gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n280_), .A2(KEYINPUT21), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  OAI211_X1 g084(.A(KEYINPUT89), .B(new_n278_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(new_n284_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT1), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G155gat), .A3(G162gat), .ZN(new_n299_));
  OR2_X1    g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n296_), .A2(new_n297_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G141gat), .ZN(new_n302_));
  INV_X1    g101(.A(G148gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT86), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT86), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(G141gat), .B2(G148gat), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n304_), .A2(new_n306_), .B1(G141gat), .B2(G148gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n300_), .A2(new_n293_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n292_), .B1(KEYINPUT29), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G228gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G22gat), .B(G50gat), .Z(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n318_), .B2(KEYINPUT29), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n301_), .A2(new_n307_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  INV_X1    g125(.A(new_n322_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n324_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G78gat), .B(G106gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT91), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n330_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n323_), .A2(new_n328_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n324_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n338_), .B2(new_n329_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n321_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n321_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n333_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT23), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G183gat), .A3(G190gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n349_), .A2(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n353_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT24), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G190gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT26), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT26), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(G190gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT92), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT26), .B(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT92), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G183gat), .ZN(new_n369_));
  INV_X1    g168(.A(G183gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT25), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n365_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT22), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G169gat), .ZN(new_n381_));
  INV_X1    g180(.A(G176gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n377_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n348_), .A2(new_n350_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n385_), .B(new_n386_), .C1(G183gat), .C2(G190gat), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n359_), .A2(new_n374_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT20), .B1(new_n388_), .B2(new_n292_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n377_), .A2(KEYINPUT24), .A3(new_n355_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n372_), .A2(KEYINPUT80), .ZN(new_n391_));
  INV_X1    g190(.A(new_n369_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n366_), .B1(new_n392_), .B2(KEYINPUT80), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n390_), .B(new_n354_), .C1(new_n391_), .C2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n383_), .A3(new_n377_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n283_), .A2(new_n286_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n347_), .B1(new_n389_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n397_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n388_), .A2(new_n292_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n347_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT20), .A4(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G8gat), .B(G36gat), .Z(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n399_), .A2(new_n408_), .A3(new_n403_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT27), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n411_), .A2(KEYINPUT27), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n361_), .A2(new_n363_), .A3(KEYINPUT92), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n416_), .A2(new_n364_), .A3(new_n372_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n395_), .B1(new_n417_), .B2(new_n358_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n397_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT98), .B(KEYINPUT20), .C1(new_n418_), .C2(new_n397_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n400_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n347_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n397_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n425_), .B(KEYINPUT20), .C1(new_n397_), .C2(new_n396_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n426_), .A2(new_n347_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n408_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT99), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n415_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n426_), .A2(new_n347_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n347_), .B2(new_n423_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n432_), .A2(KEYINPUT99), .A3(new_n408_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n345_), .B(new_n414_), .C1(new_n430_), .C2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n394_), .A2(KEYINPUT30), .A3(new_n395_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT30), .B1(new_n394_), .B2(new_n395_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n435_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n435_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n436_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT83), .B(G15gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT82), .B(G43gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G127gat), .B(G134gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G120gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT31), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n451_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n439_), .A2(new_n442_), .A3(new_n448_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n318_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n325_), .A2(new_n454_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(KEYINPUT4), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n325_), .A2(KEYINPUT4), .A3(new_n454_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n463_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G29gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G85gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n467_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n450_), .A2(new_n458_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n456_), .B1(new_n480_), .B2(new_n451_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n455_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n459_), .B(new_n479_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n434_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT99), .B1(new_n432_), .B2(new_n408_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n424_), .A2(new_n427_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n429_), .A3(new_n409_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n487_), .A3(new_n415_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n478_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n414_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n477_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n467_), .A2(KEYINPUT33), .A3(new_n468_), .A4(new_n474_), .ZN(new_n493_));
  AND4_X1   g292(.A1(new_n411_), .A2(new_n492_), .A3(new_n410_), .A4(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n308_), .A2(new_n454_), .A3(new_n317_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n325_), .A2(new_n454_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT94), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n461_), .A2(new_n498_), .A3(new_n462_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n465_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n475_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(KEYINPUT95), .A3(new_n475_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n463_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n505_), .A2(new_n506_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n507_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n404_), .B2(KEYINPUT97), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n403_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n486_), .B2(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n494_), .A2(new_n509_), .B1(new_n515_), .B2(new_n478_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n340_), .A2(new_n344_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n490_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n481_), .A2(new_n482_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n459_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n484_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G43gat), .B(G50gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n524_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529_));
  INV_X1    g328(.A(G1gat), .ZN(new_n530_));
  INV_X1    g329(.A(G8gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G8gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n527_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n525_), .A2(KEYINPUT15), .A3(new_n526_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n535_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n528_), .B(new_n535_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n537_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n538_), .A2(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT78), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G169gat), .B(G197gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n547_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT79), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n277_), .A2(new_n522_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT36), .Z(new_n559_));
  OAI211_X1 g358(.A(new_n216_), .B(new_n527_), .C1(new_n253_), .C2(new_n255_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n237_), .B2(new_n542_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n562_));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n564_), .A2(KEYINPUT35), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n561_), .A2(KEYINPUT70), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT70), .B1(new_n561_), .B2(new_n565_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n564_), .A2(KEYINPUT35), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n560_), .B(new_n570_), .C1(new_n237_), .C2(new_n542_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT71), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n543_), .A2(new_n256_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n560_), .A4(new_n570_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n559_), .B1(new_n568_), .B2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n219_), .A2(new_n224_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n231_), .B1(new_n579_), .B2(new_n250_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n236_), .B1(new_n580_), .B2(new_n234_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n542_), .B1(new_n581_), .B2(new_n216_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n560_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n565_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n561_), .A2(KEYINPUT70), .A3(new_n565_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n586_), .A2(new_n587_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n577_), .A2(KEYINPUT72), .B1(new_n578_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n559_), .ZN(new_n590_));
  OR3_X1    g389(.A1(new_n588_), .A2(KEYINPUT72), .A3(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n555_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  AOI221_X4 g391(.A(KEYINPUT73), .B1(new_n572_), .B2(new_n575_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n587_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n572_), .A2(new_n575_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n559_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT74), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT73), .B1(new_n568_), .B2(new_n576_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n559_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n588_), .A2(new_n578_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(KEYINPUT37), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n592_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G127gat), .B(G155gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n535_), .B(new_n616_), .Z(new_n617_));
  INV_X1    g416(.A(new_n247_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n617_), .B(new_n245_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT77), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n609_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n554_), .A2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n530_), .A3(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n607_), .B1(new_n599_), .B2(new_n604_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n522_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT102), .ZN(new_n639_));
  INV_X1    g438(.A(new_n277_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n626_), .A3(new_n552_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n639_), .A2(new_n479_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n636_), .B1(new_n530_), .B2(new_n642_), .ZN(G1324gat));
  NOR2_X1   g442(.A1(new_n639_), .A2(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n488_), .A2(new_n414_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n531_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n629_), .A2(new_n531_), .A3(new_n645_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT103), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n521_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n644_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT41), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n629_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n644_), .B2(new_n517_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT42), .Z(new_n661_));
  NAND3_X1  g460(.A1(new_n629_), .A2(new_n659_), .A3(new_n517_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  INV_X1    g462(.A(new_n637_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n626_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n554_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n478_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n275_), .A2(new_n627_), .A3(new_n552_), .A4(new_n276_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n603_), .B1(new_n602_), .B2(new_n559_), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT74), .B(new_n590_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n608_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n592_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(new_n522_), .A3(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n488_), .A2(new_n489_), .A3(new_n414_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n410_), .A2(new_n411_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n509_), .A2(new_n678_), .A3(new_n493_), .A4(new_n492_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n515_), .A2(new_n478_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n517_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n521_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n484_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n676_), .B1(new_n609_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n669_), .B1(new_n675_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT104), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n674_), .B2(new_n522_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n609_), .A2(new_n684_), .A3(new_n676_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n668_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n687_), .A2(new_n688_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(KEYINPUT44), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n633_), .A2(G29gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n667_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(new_n645_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n691_), .B2(KEYINPUT44), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT104), .B(new_n668_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT105), .B(new_n700_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT105), .B1(new_n694_), .B2(new_n700_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT106), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(G36gat), .A4(new_n703_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n645_), .A2(KEYINPUT107), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n645_), .A2(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n666_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n712_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n712_), .A2(KEYINPUT46), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  NAND2_X1  g523(.A1(new_n696_), .A2(new_n654_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n521_), .A2(G43gat), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n725_), .A2(G43gat), .B1(new_n666_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n666_), .B2(new_n517_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n517_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n696_), .B2(new_n730_), .ZN(G1331gat));
  INV_X1    g530(.A(new_n552_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n277_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n522_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n628_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n633_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT109), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n553_), .A2(new_n626_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n639_), .A2(new_n640_), .A3(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(G57gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n479_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n739_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n739_), .B2(new_n716_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT48), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n743_), .A3(new_n716_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n739_), .B2(new_n654_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n735_), .A2(new_n748_), .A3(new_n654_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT111), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n755_), .A3(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1334gat));
  INV_X1    g556(.A(G78gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n739_), .B2(new_n517_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n735_), .A2(new_n758_), .A3(new_n517_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n689_), .A2(new_n690_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n733_), .A2(new_n626_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n479_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n734_), .A2(new_n665_), .ZN(new_n768_));
  INV_X1    g567(.A(G85gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n633_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n768_), .B2(new_n645_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n766_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n716_), .A2(new_n202_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT113), .ZN(G1337gat));
  AOI21_X1  g575(.A(new_n221_), .B1(new_n773_), .B2(new_n654_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n654_), .A2(new_n205_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n768_), .B2(new_n778_), .ZN(new_n779_));
  XOR2_X1   g578(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n768_), .A2(new_n206_), .A3(new_n517_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n773_), .A2(new_n517_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n206_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g588(.A1(new_n521_), .A2(new_n434_), .A3(new_n632_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT119), .Z(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n544_), .A2(new_n536_), .A3(new_n546_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n551_), .B1(new_n545_), .B2(new_n537_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n547_), .A2(new_n551_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n273_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n272_), .A2(new_n552_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT55), .B1(new_n259_), .B2(new_n260_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n261_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n259_), .A2(KEYINPUT55), .A3(new_n260_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n269_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n798_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n802_), .B2(KEYINPUT118), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n797_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n792_), .B1(new_n808_), .B2(new_n637_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n798_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n800_), .A2(new_n801_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n269_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n807_), .B(new_n810_), .C1(new_n812_), .C2(KEYINPUT118), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n796_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(KEYINPUT57), .A3(new_n664_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n802_), .A2(new_n803_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n272_), .A2(new_n795_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n819_), .B2(new_n804_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n812_), .A2(KEYINPUT58), .A3(new_n817_), .A4(new_n818_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n609_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n809_), .A2(new_n815_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n627_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n738_), .B(KEYINPUT116), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT117), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n277_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n674_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(KEYINPUT54), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n828_), .A2(KEYINPUT117), .A3(new_n826_), .A4(new_n674_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n791_), .B1(new_n824_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n552_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n823_), .A2(new_n627_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n837_), .C2(new_n791_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n553_), .B(new_n842_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n836_), .B1(new_n846_), .B2(new_n835_), .ZN(G1340gat));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  AOI21_X1  g647(.A(G120gat), .B1(new_n277_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n848_), .B2(G120gat), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n834_), .B(new_n850_), .C1(new_n849_), .C2(new_n852_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n640_), .B(new_n842_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n854_));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n834_), .A2(new_n857_), .A3(new_n626_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n627_), .B(new_n842_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n857_), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n834_), .A2(new_n861_), .A3(new_n637_), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n674_), .B(new_n842_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n837_), .A2(new_n654_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n716_), .A2(new_n345_), .A3(new_n632_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n732_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n302_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n640_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n303_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n867_), .A2(new_n627_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n867_), .B2(new_n674_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n664_), .A2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n867_), .B2(new_n876_), .ZN(G1347gat));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n824_), .A2(new_n833_), .ZN(new_n879_));
  AND4_X1   g678(.A1(new_n345_), .A2(new_n716_), .A3(new_n654_), .A4(new_n632_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n732_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n882_), .B2(new_n378_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n884_));
  OAI211_X1 g683(.A(KEYINPUT62), .B(G169gat), .C1(new_n881_), .C2(new_n732_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(G1348gat));
  NOR2_X1   g685(.A1(new_n881_), .A2(new_n640_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n382_), .ZN(G1349gat));
  NAND2_X1  g687(.A1(new_n370_), .A2(KEYINPUT123), .ZN(new_n889_));
  INV_X1    g688(.A(new_n881_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n626_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n373_), .B1(KEYINPUT123), .B2(G183gat), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n881_), .A2(new_n627_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT124), .B1(new_n891_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n626_), .A3(new_n892_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n881_), .A2(new_n627_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n896_), .B(new_n897_), .C1(new_n898_), .C2(new_n889_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n881_), .B2(new_n674_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n637_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n881_), .B2(new_n902_), .ZN(G1351gat));
  NAND2_X1  g702(.A1(new_n716_), .A2(new_n489_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n837_), .A2(new_n654_), .A3(new_n732_), .A4(new_n904_), .ZN(new_n905_));
  OR3_X1    g704(.A1(new_n905_), .A2(KEYINPUT126), .A3(G197gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(KEYINPUT126), .B1(new_n905_), .B2(G197gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(G197gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT125), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n905_), .A2(new_n910_), .A3(G197gat), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n906_), .A2(new_n907_), .B1(new_n909_), .B2(new_n911_), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n837_), .A2(new_n654_), .A3(new_n904_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n277_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n914_), .B(new_n915_), .Z(G1353gat));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n626_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n917_), .B2(new_n920_), .ZN(G1354gat));
  INV_X1    g720(.A(new_n913_), .ZN(new_n922_));
  OR3_X1    g721(.A1(new_n922_), .A2(G218gat), .A3(new_n664_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G218gat), .B1(new_n922_), .B2(new_n674_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1355gat));
endmodule


