//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT3), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT2), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n206_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n209_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n211_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n204_), .B1(new_n213_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n213_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n202_), .B(new_n203_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n218_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(KEYINPUT4), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G225gat), .A2(G233gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n218_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n204_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G1gat), .B(G29gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G85gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n230_), .A2(new_n237_), .A3(new_n231_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G227gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(G15gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n244_), .B(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT79), .B(G183gat), .Z(new_n250_));
  AOI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(KEYINPUT25), .ZN(new_n251_));
  INV_X1    g050(.A(G190gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT26), .B1(new_n252_), .B2(KEYINPUT80), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(KEYINPUT26), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(KEYINPUT80), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n257_));
  INV_X1    g056(.A(G169gat), .ZN(new_n258_));
  INV_X1    g057(.A(G176gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT24), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n256_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT82), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n260_), .A2(KEYINPUT24), .A3(new_n261_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272_));
  OR3_X1    g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT22), .B(G169gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n259_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n269_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT84), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT79), .B(G183gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n252_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n280_), .A2(KEYINPUT84), .B1(new_n266_), .B2(new_n283_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n268_), .A2(new_n275_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT85), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(KEYINPUT85), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n248_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(new_n248_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n290_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n241_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n280_), .B1(new_n266_), .B2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n260_), .A2(KEYINPUT24), .A3(new_n269_), .A4(new_n261_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(KEYINPUT89), .A3(new_n304_), .A4(new_n264_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n264_), .A2(new_n304_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT89), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n298_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n311_));
  INV_X1    g110(.A(G197gat), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(G204gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(G204gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT21), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n317_), .B2(new_n314_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n317_), .B2(new_n314_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n315_), .B(new_n316_), .C1(new_n319_), .C2(KEYINPUT21), .ZN(new_n320_));
  INV_X1    g119(.A(new_n316_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(KEYINPUT21), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n310_), .A2(new_n311_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n320_), .A2(new_n322_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n285_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT90), .B1(new_n326_), .B2(new_n309_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT88), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  AOI211_X1 g132(.A(new_n325_), .B(new_n331_), .C1(new_n326_), .C2(new_n309_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n285_), .A2(new_n326_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n333_), .A2(new_n337_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n333_), .A2(KEYINPUT98), .A3(new_n337_), .A4(new_n342_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n298_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n306_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT20), .B1(new_n348_), .B2(new_n323_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n331_), .B1(new_n335_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n341_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT27), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n343_), .A2(KEYINPUT91), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n333_), .A2(new_n337_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n341_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT27), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT91), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n333_), .A2(new_n359_), .A3(new_n337_), .A4(new_n342_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .A4(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(G78gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G106gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n365_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n227_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n323_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G22gat), .B(G50gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n370_), .B(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n296_), .A2(new_n362_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT33), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n240_), .B(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n224_), .A2(new_n225_), .A3(new_n229_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n224_), .A2(KEYINPUT94), .A3(new_n225_), .A4(new_n229_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT93), .B1(new_n220_), .B2(new_n223_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n225_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n220_), .A2(KEYINPUT93), .A3(new_n223_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n237_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT95), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(KEYINPUT95), .A3(new_n389_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n380_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(new_n360_), .A3(new_n357_), .A4(new_n355_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n351_), .A2(new_n396_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT96), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n396_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n333_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n333_), .B2(new_n399_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n397_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT97), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n397_), .B(KEYINPUT97), .C1(new_n400_), .C2(new_n401_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n376_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n376_), .A2(new_n241_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n362_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n294_), .A2(new_n295_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n378_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G29gat), .B(G36gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G43gat), .B(G50gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n416_), .B(KEYINPUT78), .Z(new_n417_));
  XNOR2_X1  g216(.A(G15gat), .B(G22gat), .ZN(new_n418_));
  INV_X1    g217(.A(G1gat), .ZN(new_n419_));
  INV_X1    g218(.A(G8gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G8gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n417_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G229gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(new_n417_), .A2(new_n424_), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n430_));
  XNOR2_X1  g229(.A(new_n416_), .B(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n424_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n426_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G113gat), .B(G141gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G169gat), .B(G197gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n428_), .A2(new_n433_), .A3(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n413_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT66), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G99gat), .A2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT6), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G99gat), .A3(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G85gat), .ZN(new_n454_));
  INV_X1    g253(.A(G92gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(KEYINPUT9), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n457_), .A2(KEYINPUT9), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n449_), .A2(new_n453_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n456_), .A2(new_n457_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n446_), .A2(new_n448_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n464_));
  INV_X1    g263(.A(G99gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n451_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n462_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n449_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT8), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n462_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n461_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G57gat), .B(G64gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G71gat), .B(G78gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT11), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n478_));
  INV_X1    g277(.A(new_n476_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n475_), .A2(KEYINPUT11), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT12), .B1(new_n474_), .B2(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n471_), .A2(new_n472_), .A3(new_n462_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n472_), .B1(new_n471_), .B2(new_n462_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n460_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n487_));
  INV_X1    g286(.A(new_n482_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n482_), .B(new_n460_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT64), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT65), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n491_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n474_), .A2(new_n482_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n491_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n493_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G120gat), .B(G148gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT5), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G176gat), .B(G204gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n444_), .B1(new_n503_), .B2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n499_), .A2(KEYINPUT66), .A3(new_n502_), .A4(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n503_), .A2(new_n508_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n511_), .A2(KEYINPUT67), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT67), .B1(new_n511_), .B2(new_n512_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G134gat), .B(G162gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT73), .ZN(new_n520_));
  XOR2_X1   g319(.A(G190gat), .B(G218gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n431_), .A2(new_n486_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n474_), .A2(new_n416_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT69), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(KEYINPUT69), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n533_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n526_), .B(new_n527_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n526_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT74), .B1(new_n524_), .B2(new_n525_), .ZN(new_n546_));
  OAI221_X1 g345(.A(new_n541_), .B1(new_n535_), .B2(new_n539_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n543_), .B(new_n547_), .C1(new_n549_), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n424_), .B(KEYINPUT76), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT77), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n557_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n482_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(new_n482_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n556_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n556_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n568_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n561_), .A2(new_n562_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n571_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n518_), .A2(new_n555_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n443_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n241_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n578_), .A2(G1gat), .A3(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT38), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT38), .ZN(new_n582_));
  INV_X1    g381(.A(new_n548_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n413_), .A2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n518_), .A2(new_n442_), .A3(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G1gat), .B1(new_n586_), .B2(new_n579_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n581_), .A2(new_n582_), .A3(new_n587_), .ZN(G1324gat));
  INV_X1    g387(.A(new_n578_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n362_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n420_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594_));
  AND4_X1   g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(G8gat), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n420_), .B1(KEYINPUT99), .B2(KEYINPUT39), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n593_), .A2(new_n596_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g398(.A(G15gat), .B1(new_n586_), .B2(new_n412_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT41), .Z(new_n601_));
  NAND3_X1  g400(.A1(new_n589_), .A2(new_n246_), .A3(new_n411_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1326gat));
  OR3_X1    g402(.A1(new_n578_), .A2(G22gat), .A3(new_n376_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G22gat), .B1(new_n586_), .B2(new_n376_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n605_), .A2(KEYINPUT42), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(KEYINPUT42), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(G1327gat));
  INV_X1    g409(.A(new_n576_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n518_), .A2(new_n442_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT43), .B1(new_n413_), .B2(new_n554_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n411_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n615_), .B(new_n555_), .C1(new_n616_), .C2(new_n378_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n613_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT101), .B1(new_n618_), .B2(KEYINPUT44), .ZN(new_n619_));
  INV_X1    g418(.A(new_n617_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n406_), .A2(new_n376_), .B1(new_n362_), .B2(new_n408_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n377_), .B1(new_n621_), .B2(new_n411_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n615_), .B1(new_n622_), .B2(new_n555_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n612_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT44), .B(new_n612_), .C1(new_n620_), .C2(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G29gat), .B1(new_n630_), .B2(new_n579_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n576_), .A2(new_n583_), .A3(KEYINPUT102), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n611_), .B2(new_n548_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n518_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n622_), .A2(new_n441_), .A3(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(KEYINPUT103), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n579_), .A2(G29gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT104), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n631_), .B1(new_n639_), .B2(new_n641_), .ZN(G1328gat));
  XNOR2_X1  g441(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(G36gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n629_), .A2(new_n590_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n628_), .B2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n637_), .A2(new_n645_), .A3(new_n638_), .A4(new_n590_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT45), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n644_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n646_), .B1(new_n619_), .B2(new_n627_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n653_), .B(new_n643_), .C1(new_n645_), .C2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1329gat));
  NAND2_X1  g455(.A1(new_n411_), .A2(G43gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n629_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n657_), .B(new_n658_), .C1(new_n619_), .C2(new_n627_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n639_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G43gat), .B1(new_n660_), .B2(new_n411_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT47), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n661_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT47), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n663_), .B(new_n664_), .C1(new_n630_), .C2(new_n657_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1330gat));
  INV_X1    g465(.A(new_n376_), .ZN(new_n667_));
  INV_X1    g466(.A(G50gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT107), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n660_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n629_), .A2(new_n667_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n628_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n672_), .B1(new_n675_), .B2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n619_), .B2(new_n627_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(KEYINPUT106), .A3(new_n668_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n671_), .B1(new_n676_), .B2(new_n678_), .ZN(G1331gat));
  NAND4_X1  g478(.A1(new_n584_), .A2(new_n442_), .A3(new_n518_), .A4(new_n611_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G57gat), .B1(new_n680_), .B2(new_n579_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n622_), .A2(KEYINPUT108), .A3(new_n442_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n516_), .A2(new_n517_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT108), .B1(new_n622_), .B2(new_n442_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n576_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n579_), .A2(G57gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n681_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT109), .Z(G1332gat));
  OAI21_X1  g490(.A(G64gat), .B1(new_n680_), .B2(new_n362_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT48), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n362_), .A2(G64gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n688_), .B2(new_n694_), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n680_), .B2(new_n412_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT49), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n412_), .A2(G71gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n688_), .B2(new_n698_), .ZN(G1334gat));
  OAI21_X1  g498(.A(G78gat), .B1(new_n680_), .B2(new_n376_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT50), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n667_), .A2(new_n367_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n688_), .B2(new_n702_), .ZN(G1335gat));
  NAND2_X1  g502(.A1(new_n634_), .A2(new_n632_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n241_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n518_), .A2(new_n442_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n611_), .B(new_n706_), .C1(new_n614_), .C2(new_n617_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n241_), .A2(G85gat), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT110), .Z(new_n709_));
  AOI22_X1  g508(.A1(new_n705_), .A2(new_n454_), .B1(new_n707_), .B2(new_n709_), .ZN(G1336gat));
  NAND2_X1  g509(.A1(new_n686_), .A2(new_n704_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n455_), .B1(new_n711_), .B2(new_n362_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n712_), .A2(KEYINPUT111), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(KEYINPUT111), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n362_), .A2(new_n455_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n713_), .A2(new_n714_), .B1(new_n707_), .B2(new_n715_), .ZN(G1337gat));
  NOR2_X1   g515(.A1(new_n706_), .A2(new_n611_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n411_), .B(new_n717_), .C1(new_n620_), .C2(new_n623_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT112), .B1(new_n718_), .B2(G99gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n411_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n721_));
  OAI22_X1  g520(.A1(new_n719_), .A2(new_n720_), .B1(new_n711_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n722_), .B(new_n724_), .ZN(G1338gat));
  OAI211_X1 g524(.A(new_n667_), .B(new_n717_), .C1(new_n620_), .C2(new_n623_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G106gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G106gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n376_), .A2(G106gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n728_), .A2(new_n729_), .B1(new_n711_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g532(.A(KEYINPUT119), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(KEYINPUT59), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n687_), .A2(new_n516_), .A3(new_n442_), .A4(new_n517_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n737_), .B(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n425_), .A2(new_n426_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n429_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n438_), .A3(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n440_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n441_), .A2(new_n511_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n493_), .B1(new_n474_), .B2(new_n482_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n483_), .A2(new_n489_), .B1(new_n747_), .B2(new_n497_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(KEYINPUT55), .A3(new_n496_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT55), .B1(new_n748_), .B2(new_n496_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(KEYINPUT115), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n499_), .A2(KEYINPUT115), .A3(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n474_), .A2(KEYINPUT12), .A3(new_n482_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n487_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n491_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT116), .B1(new_n756_), .B2(new_n493_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n501_), .B1(new_n483_), .B2(new_n489_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n494_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n753_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n508_), .B1(new_n751_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n499_), .A2(new_n752_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(KEYINPUT116), .A3(new_n493_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n759_), .B1(new_n758_), .B2(new_n494_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n767_), .A2(new_n770_), .A3(new_n749_), .A4(new_n753_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n508_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n746_), .B1(new_n764_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n745_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT117), .B(new_n746_), .C1(new_n764_), .C2(new_n772_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n548_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT57), .B(new_n548_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n744_), .A2(new_n511_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n508_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(KEYINPUT118), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n764_), .A2(new_n772_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(KEYINPUT118), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n554_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n783_), .B(KEYINPUT58), .C1(new_n784_), .C2(KEYINPUT118), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(new_n780_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n740_), .B1(new_n790_), .B2(new_n576_), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n590_), .A2(new_n412_), .A3(new_n579_), .A4(new_n667_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n736_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n795_));
  AOI22_X1  g594(.A1(new_n777_), .A2(new_n778_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n611_), .B1(new_n796_), .B2(new_n780_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n792_), .B(new_n795_), .C1(new_n797_), .C2(new_n740_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n441_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G113gat), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n791_), .A2(new_n793_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n441_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT120), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(new_n806_), .A3(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1340gat));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n684_), .B2(KEYINPUT60), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n801_), .B(new_n810_), .C1(KEYINPUT60), .C2(new_n809_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n794_), .A2(new_n798_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n518_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(new_n809_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n801_), .B2(new_n611_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n611_), .A2(G127gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT121), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n812_), .B2(new_n817_), .ZN(G1342gat));
  INV_X1    g617(.A(G134gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n801_), .A2(new_n819_), .A3(new_n583_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n812_), .A2(new_n555_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n819_), .ZN(G1343gat));
  INV_X1    g621(.A(new_n791_), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n590_), .A2(new_n579_), .A3(new_n411_), .A4(new_n376_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n441_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g627(.A1(new_n825_), .A2(new_n684_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT122), .B(G148gat), .Z(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1345gat));
  XNOR2_X1  g630(.A(KEYINPUT61), .B(G155gat), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT123), .B1(new_n825_), .B2(new_n576_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n825_), .A2(KEYINPUT123), .A3(new_n576_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n836_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n834_), .A3(new_n832_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n825_), .B2(new_n554_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n548_), .A2(G162gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n825_), .B2(new_n842_), .ZN(G1347gat));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n791_), .A2(new_n362_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n376_), .A3(new_n296_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n442_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n847_), .B2(new_n258_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n276_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT62), .B(G169gat), .C1(new_n846_), .C2(new_n442_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(G1348gat));
  OAI21_X1  g650(.A(new_n518_), .B1(KEYINPUT124), .B2(G176gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n846_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(KEYINPUT124), .A2(G176gat), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT125), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n853_), .B(new_n855_), .ZN(G1349gat));
  NOR3_X1   g655(.A1(new_n846_), .A2(new_n299_), .A3(new_n576_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n846_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n611_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n282_), .B2(new_n859_), .ZN(G1350gat));
  OAI21_X1  g659(.A(G190gat), .B1(new_n846_), .B2(new_n554_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n583_), .A2(new_n300_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n846_), .B2(new_n862_), .ZN(G1351gat));
  NOR3_X1   g662(.A1(new_n411_), .A2(new_n241_), .A3(new_n376_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n845_), .A2(G197gat), .A3(new_n441_), .A4(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n865_), .A2(KEYINPUT126), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(KEYINPUT126), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n845_), .A2(new_n864_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n312_), .B1(new_n868_), .B2(new_n442_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(G1352gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n684_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT127), .B(G204gat), .Z(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1353gat));
  NOR2_X1   g672(.A1(new_n868_), .A2(new_n576_), .ZN(new_n874_));
  OR2_X1    g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT63), .B(G211gat), .Z(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n874_), .B2(new_n877_), .ZN(G1354gat));
  OAI21_X1  g677(.A(G218gat), .B1(new_n868_), .B2(new_n554_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n548_), .A2(G218gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n868_), .B2(new_n880_), .ZN(G1355gat));
endmodule


