//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(KEYINPUT69), .ZN(new_n204_));
  XOR2_X1   g003(.A(G43gat), .B(G50gat), .Z(new_n205_));
  OR3_X1    g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n205_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT7), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n215_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n215_), .B(new_n226_), .C1(new_n218_), .C2(new_n224_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n221_), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n213_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n239_), .B(KEYINPUT34), .Z(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT68), .B(KEYINPUT35), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n210_), .A2(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n237_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT65), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n242_), .B1(new_n208_), .B2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n240_), .A2(new_n241_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT36), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G190gat), .B(G218gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT71), .ZN(new_n256_));
  XOR2_X1   g055(.A(G134gat), .B(G162gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(KEYINPUT36), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT37), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT37), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n264_), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G127gat), .B(G155gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT16), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G183gat), .B(G211gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT17), .ZN(new_n271_));
  XOR2_X1   g070(.A(G71gat), .B(G78gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(G57gat), .B(G64gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(KEYINPUT11), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT66), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n272_), .B(new_n276_), .C1(KEYINPUT11), .C2(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(KEYINPUT11), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G15gat), .B(G22gat), .ZN(new_n281_));
  INV_X1    g080(.A(G1gat), .ZN(new_n282_));
  INV_X1    g081(.A(G8gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT14), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G1gat), .B(G8gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G231gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n280_), .B(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n271_), .B1(new_n290_), .B2(KEYINPUT73), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(KEYINPUT73), .B2(new_n290_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n270_), .A2(KEYINPUT17), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT72), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n266_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT74), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n248_), .B2(new_n280_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n278_), .A2(new_n279_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n275_), .A2(new_n277_), .B1(KEYINPUT11), .B2(new_n273_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n244_), .A2(new_n302_), .A3(new_n247_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n280_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n299_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G230gat), .A2(G233gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n303_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n302_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G120gat), .B(G148gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n308_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n308_), .B2(new_n312_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT13), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(KEYINPUT13), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n298_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT96), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  OR2_X1    g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n329_), .A2(KEYINPUT21), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G197gat), .A2(G204gat), .ZN(new_n336_));
  AND2_X1   g135(.A1(G197gat), .A2(G204gat), .ZN(new_n337_));
  AND2_X1   g136(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n339_));
  OAI22_X1  g138(.A1(new_n336_), .A2(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n334_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n341_));
  OAI221_X1 g140(.A(KEYINPUT84), .B1(new_n337_), .B2(new_n336_), .C1(new_n339_), .C2(new_n338_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n333_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT23), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(G183gat), .A3(G190gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n345_), .A2(new_n347_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(G169gat), .B2(G176gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n349_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355_));
  INV_X1    g154(.A(G183gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(KEYINPUT25), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(G190gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT25), .B(G183gat), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n357_), .B(new_n358_), .C1(new_n359_), .C2(new_n355_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n344_), .A2(new_n346_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n362_));
  INV_X1    g161(.A(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G176gat), .ZN(new_n368_));
  INV_X1    g167(.A(G169gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT79), .B1(new_n369_), .B2(KEYINPUT22), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT22), .B(G169gat), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n368_), .B(new_n370_), .C1(new_n371_), .C2(KEYINPUT79), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n354_), .A2(new_n360_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n328_), .B1(new_n343_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT19), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT88), .Z(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n368_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n359_), .A2(new_n358_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n381_));
  AOI221_X4 g180(.A(KEYINPUT89), .B1(new_n349_), .B2(new_n348_), .C1(new_n345_), .C2(new_n347_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT89), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n345_), .A2(new_n347_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n349_), .A2(new_n348_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n381_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT90), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT90), .B(new_n381_), .C1(new_n382_), .C2(new_n386_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n380_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n374_), .B(new_n377_), .C1(new_n391_), .C2(new_n343_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT20), .B1(new_n343_), .B2(new_n373_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n340_), .A2(new_n335_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n394_), .A2(new_n342_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n333_), .ZN(new_n396_));
  AND4_X1   g195(.A1(new_n395_), .A2(new_n387_), .A3(new_n396_), .A4(new_n379_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n376_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n384_), .A2(new_n385_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT89), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n350_), .A2(new_n383_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT90), .B1(new_n410_), .B2(new_n381_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n390_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n343_), .B(new_n379_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n376_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n395_), .A2(new_n396_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n367_), .A2(new_n372_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n360_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n328_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT20), .B1(new_n415_), .B2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n379_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n415_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n404_), .B(new_n420_), .C1(new_n423_), .C2(new_n377_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n406_), .A2(KEYINPUT27), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT95), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT95), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n406_), .A2(new_n424_), .A3(new_n427_), .A4(KEYINPUT27), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n374_), .B1(new_n391_), .B2(new_n343_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n377_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(KEYINPUT92), .A3(new_n404_), .A4(new_n420_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n420_), .B1(new_n423_), .B2(new_n377_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n405_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n429_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT0), .B(G57gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT80), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G127gat), .B(G134gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G120gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n449_), .B(new_n451_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n448_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT2), .ZN(new_n456_));
  INV_X1    g255(.A(G141gat), .ZN(new_n457_));
  INV_X1    g256(.A(G148gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT3), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n459_), .A2(new_n461_), .A3(new_n462_), .A4(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G141gat), .B(G148gat), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(KEYINPUT1), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n465_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n466_), .A2(KEYINPUT1), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT4), .B1(new_n455_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n455_), .A2(new_n474_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n454_), .A2(new_n473_), .A3(new_n468_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI211_X1 g277(.A(new_n447_), .B(new_n475_), .C1(new_n478_), .C2(KEYINPUT4), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n447_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n446_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(KEYINPUT4), .ZN(new_n483_));
  INV_X1    g282(.A(new_n447_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n475_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n445_), .A3(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n482_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT81), .B(KEYINPUT28), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n474_), .A2(KEYINPUT29), .ZN(new_n492_));
  XOR2_X1   g291(.A(G22gat), .B(G50gat), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n492_), .A2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n491_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(KEYINPUT82), .A2(G233gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(KEYINPUT82), .A2(G233gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(G228gat), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n415_), .B2(KEYINPUT85), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n474_), .A2(KEYINPUT29), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n415_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n415_), .B(new_n506_), .C1(KEYINPUT85), .C2(new_n504_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G78gat), .B(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n508_), .A2(KEYINPUT86), .A3(new_n509_), .A4(new_n511_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n508_), .A2(new_n509_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n510_), .ZN(new_n519_));
  AOI211_X1 g318(.A(KEYINPUT87), .B(new_n511_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n501_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n510_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n501_), .A2(new_n523_), .A3(new_n512_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n489_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n327_), .B1(new_n441_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(KEYINPUT87), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n518_), .A2(new_n517_), .A3(new_n510_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n501_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n524_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n488_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n533_), .A2(KEYINPUT96), .A3(new_n440_), .A4(new_n429_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n399_), .A2(KEYINPUT32), .A3(new_n404_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT94), .Z(new_n537_));
  OAI211_X1 g336(.A(new_n488_), .B(new_n535_), .C1(new_n436_), .C2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT33), .B(new_n446_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT93), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n484_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n445_), .B1(new_n478_), .B2(new_n447_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT33), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n482_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n445_), .B1(new_n486_), .B2(new_n480_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT33), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n538_), .B1(new_n548_), .B2(new_n438_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n524_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n526_), .A2(new_n534_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G227gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(G15gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT30), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n418_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(new_n455_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G71gat), .B(G99gat), .ZN(new_n559_));
  INV_X1    g358(.A(G43gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT31), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n429_), .A2(new_n550_), .A3(new_n440_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT97), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n429_), .A2(new_n550_), .A3(new_n440_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n489_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n552_), .A2(new_n566_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT75), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n208_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n287_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n210_), .A2(new_n287_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n578_), .A2(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G113gat), .B(G141gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n574_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n326_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n282_), .B1(KEYINPUT98), .B2(KEYINPUT38), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n594_), .A2(new_n489_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(KEYINPUT98), .A2(KEYINPUT38), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n262_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n574_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n325_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n600_), .A2(new_n591_), .A3(new_n601_), .A4(new_n296_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT99), .Z(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n603_), .B2(new_n489_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(new_n441_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G8gat), .B1(new_n602_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT39), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n441_), .A2(new_n283_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n594_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  NOR2_X1   g410(.A1(new_n603_), .A2(new_n566_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n612_), .A2(KEYINPUT41), .A3(new_n554_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT41), .B1(new_n612_), .B2(new_n554_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n565_), .A2(new_n554_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n594_), .A2(KEYINPUT100), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT100), .B1(new_n594_), .B2(new_n615_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .A4(new_n617_), .ZN(G1326gat));
  NAND2_X1  g417(.A1(new_n531_), .A2(new_n532_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT101), .ZN(new_n620_));
  OAI21_X1  g419(.A(G22gat), .B1(new_n603_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT42), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(G22gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT102), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n622_), .B1(new_n594_), .B2(new_n624_), .ZN(G1327gat));
  INV_X1    g424(.A(KEYINPUT104), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT44), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n325_), .A2(new_n592_), .A3(new_n296_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT43), .B1(new_n574_), .B2(new_n266_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n266_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n619_), .A2(new_n429_), .A3(new_n489_), .A4(new_n440_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n633_), .A2(new_n327_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n565_), .B1(new_n634_), .B2(new_n534_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n572_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n631_), .B(new_n632_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n629_), .B1(new_n630_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n627_), .B1(new_n638_), .B2(KEYINPUT103), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n640_), .B(new_n629_), .C1(new_n630_), .C2(new_n637_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n626_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n552_), .A2(new_n566_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n636_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n632_), .B1(new_n645_), .B2(new_n631_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n574_), .A2(KEYINPUT43), .A3(new_n266_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n628_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n640_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n638_), .A2(KEYINPUT103), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(KEYINPUT104), .A3(new_n627_), .A4(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n642_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n638_), .A2(KEYINPUT44), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(G29gat), .A3(new_n488_), .A4(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n262_), .A2(new_n296_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n593_), .A2(new_n601_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n488_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n654_), .A2(KEYINPUT105), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1328gat));
  XNOR2_X1  g463(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(G36gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n653_), .A2(new_n441_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n652_), .B2(new_n669_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n656_), .A2(G36gat), .A3(new_n606_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n666_), .B1(new_n670_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n668_), .B1(new_n642_), .B2(new_n651_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n673_), .B(new_n665_), .C1(new_n676_), .C2(new_n667_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1329gat));
  NAND4_X1  g477(.A1(new_n652_), .A2(G43gat), .A3(new_n565_), .A4(new_n653_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G43gat), .B1(new_n657_), .B2(new_n565_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT47), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n679_), .A2(new_n684_), .A3(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1330gat));
  NAND4_X1  g485(.A1(new_n652_), .A2(G50gat), .A3(new_n619_), .A4(new_n653_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n620_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G50gat), .B1(new_n657_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n687_), .A2(KEYINPUT108), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1331gat));
  NOR4_X1   g494(.A1(new_n298_), .A2(new_n574_), .A3(new_n591_), .A4(new_n601_), .ZN(new_n696_));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n488_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n296_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n591_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n600_), .A2(new_n325_), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n489_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(G1332gat));
  OAI21_X1  g502(.A(G64gat), .B1(new_n701_), .B2(new_n606_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n696_), .A2(new_n707_), .A3(new_n441_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n701_), .B2(new_n566_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n696_), .A2(new_n713_), .A3(new_n565_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1334gat));
  OAI21_X1  g514(.A(G78gat), .B1(new_n701_), .B2(new_n620_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G78gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n696_), .A2(new_n719_), .A3(new_n688_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1335gat));
  NAND4_X1  g520(.A1(new_n645_), .A2(new_n592_), .A3(new_n325_), .A4(new_n655_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n211_), .A3(new_n488_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n325_), .A2(new_n592_), .A3(new_n699_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n630_), .B2(new_n637_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(new_n488_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(new_n211_), .ZN(G1336gat));
  NAND3_X1  g527(.A1(new_n723_), .A2(new_n212_), .A3(new_n441_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n726_), .A2(new_n441_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n212_), .ZN(G1337gat));
  NAND4_X1  g530(.A1(new_n723_), .A2(new_n565_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT112), .Z(new_n733_));
  AOI21_X1  g532(.A(new_n220_), .B1(new_n726_), .B2(new_n565_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n723_), .A2(new_n221_), .A3(new_n619_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n726_), .A2(new_n619_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G106gat), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT52), .B(new_n221_), .C1(new_n726_), .C2(new_n619_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g542(.A(new_n588_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n576_), .A2(new_n577_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n581_), .A2(new_n745_), .A3(new_n580_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n590_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n319_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT55), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n303_), .B(new_n304_), .C1(new_n311_), .C2(KEYINPUT12), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n309_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n309_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n303_), .A2(new_n304_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n246_), .A2(KEYINPUT65), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n243_), .B(new_n245_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n280_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT12), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n756_), .A2(new_n761_), .A3(KEYINPUT55), .A4(new_n307_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n306_), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n307_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n755_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n750_), .B1(new_n766_), .B2(new_n318_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n764_), .A2(new_n765_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n307_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n308_), .B2(new_n751_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n318_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n749_), .B1(new_n767_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n773_), .A2(KEYINPUT116), .A3(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n748_), .A2(new_n319_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n768_), .A2(new_n770_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n317_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n750_), .B(new_n318_), .C1(new_n768_), .C2(new_n770_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT58), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n631_), .B1(new_n775_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  INV_X1    g585(.A(new_n748_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(new_n322_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n771_), .B2(KEYINPUT56), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT115), .B(new_n750_), .C1(new_n766_), .C2(new_n318_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n772_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n592_), .A2(new_n320_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n786_), .B1(new_n794_), .B2(new_n599_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n792_), .A2(new_n793_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT57), .B(new_n262_), .C1(new_n796_), .C2(new_n788_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n774_), .B1(new_n773_), .B2(KEYINPUT116), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(KEYINPUT117), .A3(new_n631_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n785_), .A2(new_n795_), .A3(new_n797_), .A4(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n699_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n700_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n601_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT113), .ZN(new_n808_));
  INV_X1    g607(.A(new_n805_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT54), .B1(new_n809_), .B2(new_n325_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n805_), .A2(new_n601_), .A3(new_n811_), .A4(new_n806_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n803_), .A2(new_n813_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n489_), .B(new_n566_), .C1(new_n568_), .C2(new_n570_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n797_), .A2(new_n795_), .A3(new_n783_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n699_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n813_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n815_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n591_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G113gat), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n816_), .A2(G113gat), .A3(new_n592_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1340gat));
  NAND3_X1  g625(.A1(new_n817_), .A2(new_n325_), .A3(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G120gat), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT60), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(G120gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(G120gat), .B1(new_n325_), .B2(new_n829_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n816_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(G1341gat));
  AND2_X1   g632(.A1(new_n817_), .A2(new_n822_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n296_), .A2(G127gat), .ZN(new_n835_));
  XOR2_X1   g634(.A(new_n835_), .B(KEYINPUT119), .Z(new_n836_));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n814_), .A2(new_n296_), .A3(new_n815_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n834_), .A2(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(G1342gat));
  NAND3_X1  g638(.A1(new_n817_), .A2(new_n631_), .A3(new_n822_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G134gat), .ZN(new_n841_));
  OR3_X1    g640(.A1(new_n816_), .A2(G134gat), .A3(new_n262_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1343gat));
  NOR3_X1   g642(.A1(new_n441_), .A2(new_n489_), .A3(new_n550_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT117), .B1(new_n800_), .B2(new_n631_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n784_), .B(new_n266_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n797_), .A2(new_n795_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n296_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n813_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n566_), .B(new_n844_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n592_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT120), .B(G141gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1344gat));
  NOR2_X1   g653(.A1(new_n851_), .A2(new_n601_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n458_), .ZN(G1345gat));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n850_), .B1(new_n802_), .B2(new_n699_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n844_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n565_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n859_), .B1(new_n862_), .B2(new_n296_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n851_), .A2(KEYINPUT121), .A3(new_n699_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n858_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n859_), .A3(new_n296_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT121), .B1(new_n851_), .B2(new_n699_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n857_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n868_), .ZN(G1346gat));
  OR3_X1    g668(.A1(new_n851_), .A2(G162gat), .A3(new_n262_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G162gat), .B1(new_n851_), .B2(new_n266_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1347gat));
  NAND2_X1  g671(.A1(new_n820_), .A2(new_n620_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n606_), .A2(new_n572_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n591_), .A2(new_n371_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT122), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n820_), .A2(new_n591_), .A3(new_n620_), .A4(new_n874_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(G169gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1348gat));
  AOI21_X1  g683(.A(G176gat), .B1(new_n876_), .B2(new_n325_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n860_), .A2(new_n619_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n601_), .A2(new_n368_), .A3(new_n875_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  NOR2_X1   g687(.A1(new_n875_), .A2(new_n699_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n873_), .A2(new_n359_), .A3(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n860_), .A2(new_n619_), .A3(new_n890_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G183gat), .B1(new_n892_), .B2(new_n893_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n891_), .B1(new_n894_), .B2(new_n895_), .ZN(G1350gat));
  AND2_X1   g695(.A1(new_n599_), .A2(new_n358_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n820_), .A2(new_n620_), .A3(new_n874_), .A4(new_n897_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n873_), .A2(new_n266_), .A3(new_n875_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n363_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n898_), .C1(new_n899_), .C2(new_n363_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1351gat));
  NOR4_X1   g703(.A1(new_n860_), .A2(new_n565_), .A3(new_n525_), .A4(new_n606_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n905_), .A2(new_n906_), .A3(G197gat), .A4(new_n591_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n606_), .A2(new_n525_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n814_), .A2(new_n566_), .A3(new_n591_), .A4(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(G197gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT125), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n910_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n907_), .A2(new_n911_), .A3(new_n912_), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n905_), .A2(new_n325_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n814_), .A2(new_n566_), .A3(new_n908_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n296_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT126), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n919_), .B(new_n921_), .ZN(G1354gat));
  OR3_X1    g721(.A1(new_n916_), .A2(G218gat), .A3(new_n262_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G218gat), .B1(new_n916_), .B2(new_n266_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1355gat));
endmodule


