//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n208_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT25), .B(G183gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT26), .B1(new_n208_), .B2(KEYINPUT82), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n213_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n203_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n207_), .B1(new_n212_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n219_), .A2(new_n212_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT83), .A3(new_n207_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT30), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(KEYINPUT30), .A3(new_n224_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT84), .B(G43gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(G15gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G71gat), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n229_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n231_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  MUX2_X1   g042(.A(new_n242_), .B(new_n243_), .S(KEYINPUT85), .Z(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT31), .Z(new_n245_));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n237_), .B1(new_n231_), .B2(new_n238_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n239_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n245_), .B(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n250_), .B1(new_n239_), .B2(new_n248_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G1gat), .B(G29gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G85gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n253_), .B(new_n254_), .Z(new_n255_));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256_));
  XOR2_X1   g055(.A(G155gat), .B(G162gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT2), .ZN(new_n259_));
  OR2_X1    g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n260_), .B2(KEYINPUT87), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n260_), .A2(KEYINPUT87), .A3(KEYINPUT3), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n257_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n260_), .A4(new_n258_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n244_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n242_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n256_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n270_), .A2(KEYINPUT4), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n274_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n255_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n271_), .A2(new_n272_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT4), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n255_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n278_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n286_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n249_), .A2(new_n251_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n264_), .A2(new_n268_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n289_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT28), .B1(new_n289_), .B2(KEYINPUT29), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G22gat), .B(G50gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G78gat), .B(G106gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT90), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n304_), .A2(new_n300_), .A3(new_n305_), .A4(KEYINPUT21), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT89), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n289_), .A2(KEYINPUT29), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT88), .ZN(new_n313_));
  INV_X1    g112(.A(G228gat), .ZN(new_n314_));
  INV_X1    g113(.A(G233gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n313_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n299_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n318_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n325_));
  OAI22_X1  g124(.A1(new_n324_), .A2(new_n325_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n313_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n298_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT92), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT92), .A4(new_n298_), .ZN(new_n331_));
  OAI211_X1 g130(.A(KEYINPUT91), .B(new_n299_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n323_), .A2(new_n330_), .A3(new_n331_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n296_), .A2(new_n321_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n328_), .A2(new_n335_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n297_), .A2(new_n333_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n307_), .A2(new_n309_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT95), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n207_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n204_), .A2(KEYINPUT95), .A3(new_n206_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n210_), .A2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n347_), .A2(KEYINPUT94), .A3(new_n218_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT94), .B1(new_n347_), .B2(new_n218_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n203_), .A2(new_n215_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n341_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(KEYINPUT20), .C1(new_n225_), .C2(new_n341_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT19), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT20), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n345_), .A2(new_n351_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n341_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n225_), .A2(new_n341_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n353_), .A2(new_n355_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NOR2_X1   g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n353_), .A2(new_n355_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n362_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n370_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n340_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n340_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n375_));
  INV_X1    g174(.A(new_n368_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n353_), .A2(new_n355_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n355_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n307_), .A2(new_n309_), .A3(new_n207_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n351_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n356_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n378_), .B1(new_n362_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n376_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n374_), .A2(new_n375_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n373_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n375_), .B1(new_n374_), .B2(new_n383_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n288_), .A2(new_n339_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n333_), .A2(new_n297_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n337_), .A2(new_n338_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n279_), .A2(new_n286_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n387_), .A3(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT32), .B(new_n368_), .C1(new_n377_), .C2(new_n382_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n363_), .B1(new_n396_), .B2(new_n376_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n287_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n279_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT33), .B(new_n255_), .C1(new_n276_), .C2(new_n278_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n369_), .A2(new_n372_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n274_), .B1(new_n280_), .B2(KEYINPUT97), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(KEYINPUT97), .B2(new_n280_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n274_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n284_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n398_), .B1(new_n402_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n339_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n394_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n249_), .A2(new_n251_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n389_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G29gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT76), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G43gat), .B(G50gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT76), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n415_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT15), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G22gat), .ZN(new_n426_));
  INV_X1    g225(.A(G1gat), .ZN(new_n427_));
  INV_X1    g226(.A(G8gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT14), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G1gat), .B(G8gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n423_), .A2(new_n432_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G229gat), .A2(G233gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n423_), .B(new_n432_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G113gat), .B(G141gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G169gat), .B(G197gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n441_), .B(new_n442_), .Z(new_n443_));
  OR2_X1    g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n443_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT81), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n414_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G78gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G64gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G57gat), .ZN(new_n456_));
  INV_X1    g255(.A(G57gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G64gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n458_), .A3(KEYINPUT11), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT70), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT70), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n456_), .A2(new_n458_), .A3(new_n462_), .A4(KEYINPUT11), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n454_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n462_), .B1(new_n450_), .B2(KEYINPUT11), .ZN(new_n467_));
  INV_X1    g266(.A(new_n463_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT69), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n453_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT6), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G99gat), .A3(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT68), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n477_), .A2(new_n478_), .A3(new_n480_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  INV_X1    g283(.A(G92gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(KEYINPUT8), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT66), .B(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT65), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n492_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n491_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n500_));
  NOR2_X1   g299(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n486_), .B(new_n487_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n487_), .A2(KEYINPUT9), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n477_), .A3(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT8), .B1(new_n483_), .B2(new_n488_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n490_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n449_), .B1(new_n472_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT72), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n475_), .B1(G99gat), .B2(G106gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n478_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n480_), .A2(new_n482_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n488_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n502_), .A2(new_n477_), .A3(new_n503_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n491_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT65), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n497_), .B1(new_n496_), .B2(new_n492_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n489_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(new_n471_), .A3(new_n466_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT72), .A3(new_n449_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n524_), .A2(KEYINPUT12), .A3(new_n471_), .A4(new_n466_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT71), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n469_), .A2(new_n453_), .A3(new_n470_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n453_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT12), .A4(new_n524_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n510_), .A2(new_n526_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n524_), .B1(new_n471_), .B2(new_n466_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G230gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT64), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT73), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n472_), .A2(new_n507_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n525_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n537_), .B1(new_n545_), .B2(new_n535_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G120gat), .B(G148gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(G176gat), .B(G204gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n547_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n544_), .A2(new_n546_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n552_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(KEYINPUT75), .A3(new_n556_), .ZN(new_n557_));
  OR3_X1    g356(.A1(new_n547_), .A2(KEYINPUT75), .A3(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT13), .B1(new_n557_), .B2(new_n558_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n425_), .A2(new_n524_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT35), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n507_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n564_), .A2(new_n565_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n569_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n564_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n570_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n564_), .B2(KEYINPUT77), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT36), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n577_), .A2(KEYINPUT78), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT78), .B1(new_n577_), .B2(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n432_), .B(KEYINPUT79), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n531_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n593_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT80), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n593_), .A2(KEYINPUT80), .A3(new_n599_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n602_), .A2(new_n603_), .B1(new_n592_), .B2(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(KEYINPUT37), .B(new_n582_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n588_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n448_), .A2(new_n563_), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n427_), .A3(new_n287_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT99), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n610_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT103), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n563_), .A2(new_n605_), .A3(new_n446_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n287_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n616_), .A2(new_n387_), .B1(new_n409_), .B2(new_n339_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n388_), .B1(new_n617_), .B2(new_n412_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n586_), .B(KEYINPUT100), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT101), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n287_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G1gat), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT102), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(KEYINPUT102), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n612_), .B(new_n614_), .C1(new_n629_), .C2(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n387_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n428_), .B1(new_n622_), .B2(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT39), .Z(new_n634_));
  NAND3_X1  g433(.A1(new_n608_), .A2(new_n428_), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g436(.A1(new_n608_), .A2(new_n233_), .A3(new_n412_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n626_), .A2(new_n412_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(new_n639_), .B2(G15gat), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641_));
  AOI211_X1 g440(.A(new_n641_), .B(new_n233_), .C1(new_n626_), .C2(new_n412_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(G1326gat));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n626_), .B2(new_n392_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n608_), .A2(new_n646_), .A3(new_n392_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(G29gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n588_), .A2(new_n606_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n414_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n412_), .B1(new_n394_), .B2(new_n410_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n655_), .B(new_n652_), .C1(new_n656_), .C2(new_n389_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n605_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n563_), .A2(new_n659_), .A3(new_n446_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n663_), .B(new_n660_), .C1(new_n654_), .C2(new_n657_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n651_), .B1(new_n665_), .B2(new_n287_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n561_), .A2(new_n562_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n620_), .A2(new_n667_), .A3(new_n605_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n448_), .A2(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(G29gat), .A3(new_n393_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n666_), .A2(new_n670_), .ZN(G1328gat));
  NOR2_X1   g470(.A1(new_n387_), .A2(G36gat), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT106), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n448_), .A2(new_n668_), .A3(new_n675_), .A4(new_n672_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n674_), .A2(KEYINPUT45), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT45), .B1(new_n674_), .B2(new_n676_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n665_), .B2(new_n632_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n657_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n655_), .B1(new_n618_), .B2(new_n652_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n661_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n663_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n661_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n685_), .A2(new_n680_), .A3(new_n686_), .A4(new_n632_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G36gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n679_), .B1(new_n681_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n689_), .A2(new_n690_), .A3(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n685_), .A2(new_n632_), .A3(new_n686_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT105), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(G36gat), .A3(new_n687_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n697_), .A2(new_n691_), .A3(new_n692_), .A4(new_n679_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n694_), .A2(new_n698_), .ZN(G1329gat));
  NOR3_X1   g498(.A1(new_n669_), .A2(G43gat), .A3(new_n413_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n665_), .A2(new_n412_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(G43gat), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g502(.A(new_n669_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G50gat), .B1(new_n704_), .B2(new_n392_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n392_), .A2(G50gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n665_), .B2(new_n706_), .ZN(G1331gat));
  NOR2_X1   g506(.A1(new_n563_), .A2(new_n659_), .ZN(new_n708_));
  AND4_X1   g507(.A1(new_n618_), .A2(new_n708_), .A3(new_n620_), .A4(new_n447_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT109), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n287_), .A2(G57gat), .ZN(new_n711_));
  OR3_X1    g510(.A1(new_n710_), .A2(KEYINPUT110), .A3(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n563_), .A2(new_n659_), .A3(new_n652_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n414_), .A2(new_n446_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n457_), .B1(new_n717_), .B2(new_n393_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT110), .B1(new_n710_), .B2(new_n711_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n712_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT111), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n712_), .A2(new_n722_), .A3(new_n718_), .A4(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(new_n717_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n455_), .A3(new_n632_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n710_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n632_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(G64gat), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  OR3_X1    g531(.A1(new_n717_), .A2(G71gat), .A3(new_n413_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n727_), .A2(new_n412_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G71gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G71gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n725_), .A2(new_n739_), .A3(new_n392_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n727_), .A2(new_n392_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G78gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT50), .B(new_n739_), .C1(new_n727_), .C2(new_n392_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  NAND4_X1  g544(.A1(new_n715_), .A2(new_n619_), .A3(new_n659_), .A4(new_n667_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n484_), .A3(new_n287_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n682_), .A2(new_n683_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n446_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n667_), .A2(new_n659_), .A3(new_n750_), .ZN(new_n751_));
  OR3_X1    g550(.A1(new_n749_), .A2(KEYINPUT113), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n749_), .B2(new_n751_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(KEYINPUT114), .A3(new_n753_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n393_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n748_), .B1(new_n758_), .B2(new_n484_), .ZN(G1336gat));
  NAND3_X1  g558(.A1(new_n747_), .A2(new_n485_), .A3(new_n632_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n387_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n485_), .ZN(G1337gat));
  OAI211_X1 g561(.A(new_n747_), .B(new_n412_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n413_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n236_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n747_), .A2(new_n392_), .A3(new_n519_), .ZN(new_n767_));
  OR3_X1    g566(.A1(new_n749_), .A2(new_n339_), .A3(new_n751_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G106gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G106gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n772_), .B(new_n774_), .ZN(G1339gat));
  OAI211_X1 g574(.A(new_n607_), .B(new_n447_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT54), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n433_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n443_), .B1(new_n437_), .B2(new_n435_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n440_), .A2(new_n443_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n557_), .A2(new_n558_), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n510_), .A2(new_n526_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n533_), .A2(new_n528_), .ZN(new_n784_));
  AND4_X1   g583(.A1(KEYINPUT55), .A2(new_n543_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT55), .B1(new_n534_), .B2(new_n543_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT72), .B1(new_n525_), .B2(new_n449_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n525_), .A2(KEYINPUT72), .A3(new_n449_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n784_), .B(new_n539_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT116), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n534_), .A2(new_n792_), .A3(new_n539_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n793_), .A3(new_n537_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n552_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n797_), .B(new_n553_), .C1(new_n787_), .C2(new_n794_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n796_), .A2(new_n798_), .A3(KEYINPUT117), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n791_), .A2(new_n537_), .A3(new_n793_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n544_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n534_), .A2(KEYINPUT55), .A3(new_n543_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n552_), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT117), .A3(new_n797_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n446_), .A2(new_n554_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n782_), .B1(new_n799_), .B2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT57), .A3(new_n620_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n797_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n807_), .B1(new_n796_), .B2(KEYINPUT117), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n781_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n812_), .B1(new_n818_), .B2(new_n619_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n813_), .A2(new_n815_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n554_), .A2(new_n780_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n821_), .B(KEYINPUT58), .C1(new_n796_), .C2(new_n798_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n652_), .A3(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n811_), .A2(new_n819_), .A3(new_n826_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n827_), .A2(KEYINPUT118), .A3(new_n659_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT118), .B1(new_n827_), .B2(new_n659_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n777_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n632_), .A2(new_n392_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n413_), .A2(new_n393_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  INV_X1    g633(.A(new_n833_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n825_), .A2(new_n652_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n820_), .B2(new_n821_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n810_), .A2(new_n620_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n812_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n605_), .B1(new_n840_), .B2(new_n811_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n776_), .B(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n835_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n830_), .A2(new_n834_), .B1(new_n844_), .B2(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846_), .B2(new_n447_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n750_), .A2(G113gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n844_), .B2(new_n848_), .ZN(G1340gat));
  XNOR2_X1  g648(.A(KEYINPUT119), .B(G120gat), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n846_), .B2(new_n563_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n563_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(KEYINPUT60), .B2(new_n850_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n844_), .B2(new_n854_), .ZN(G1341gat));
  OAI21_X1  g654(.A(G127gat), .B1(new_n846_), .B2(new_n659_), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n659_), .A2(G127gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n844_), .B2(new_n857_), .ZN(G1342gat));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n845_), .B2(new_n652_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n844_), .A2(G134gat), .A3(new_n620_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n843_), .B1(new_n659_), .B2(new_n827_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n864_), .B2(new_n833_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n829_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n827_), .A2(KEYINPUT118), .A3(new_n659_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n843_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n834_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n865_), .B(new_n652_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G134gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n862_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(KEYINPUT120), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n863_), .A2(new_n873_), .ZN(G1343gat));
  NAND2_X1  g673(.A1(new_n827_), .A2(new_n659_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n777_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n632_), .A2(new_n339_), .A3(new_n393_), .A4(new_n412_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n446_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n667_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g682(.A1(new_n878_), .A2(new_n659_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT61), .B(G155gat), .Z(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  OR3_X1    g685(.A1(new_n878_), .A2(G162gat), .A3(new_n620_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G162gat), .B1(new_n878_), .B2(new_n653_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1347gat));
  INV_X1    g688(.A(G169gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n632_), .A2(new_n288_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n392_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n750_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n890_), .B1(new_n830_), .B2(new_n894_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n895_), .A2(KEYINPUT122), .A3(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT22), .B(G169gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n830_), .A2(new_n894_), .A3(new_n899_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n895_), .A2(KEYINPUT122), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n895_), .B2(KEYINPUT122), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n898_), .B(new_n900_), .C1(new_n901_), .C2(new_n902_), .ZN(G1348gat));
  NAND2_X1  g702(.A1(new_n876_), .A2(new_n339_), .ZN(new_n904_));
  INV_X1    g703(.A(G176gat), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n563_), .A4(new_n891_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n830_), .A2(new_n892_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n907_), .B2(new_n563_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT123), .B(new_n905_), .C1(new_n907_), .C2(new_n563_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n906_), .B1(new_n910_), .B2(new_n911_), .ZN(G1349gat));
  OR2_X1    g711(.A1(new_n659_), .A2(new_n210_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n907_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(KEYINPUT124), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n891_), .A2(new_n659_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n876_), .A2(new_n339_), .A3(new_n916_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n918_), .A2(new_n919_), .A3(G183gat), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n907_), .A2(new_n921_), .A3(new_n913_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n915_), .A2(new_n920_), .A3(new_n922_), .ZN(G1350gat));
  OAI21_X1  g722(.A(G190gat), .B1(new_n907_), .B2(new_n653_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n619_), .A2(new_n346_), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT126), .Z(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n907_), .B2(new_n926_), .ZN(G1351gat));
  AND3_X1   g726(.A1(new_n632_), .A2(new_n616_), .A3(new_n413_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n876_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n446_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n667_), .ZN(new_n933_));
  INV_X1    g732(.A(G204gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(KEYINPUT127), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n933_), .B(new_n935_), .ZN(G1353gat));
  NAND2_X1  g735(.A1(new_n930_), .A2(new_n605_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  AND2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(new_n937_), .B2(new_n938_), .ZN(G1354gat));
  OR3_X1    g740(.A1(new_n929_), .A2(G218gat), .A3(new_n620_), .ZN(new_n942_));
  OAI21_X1  g741(.A(G218gat), .B1(new_n929_), .B2(new_n653_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1355gat));
endmodule


