//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G71gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G43gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT79), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n206_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT76), .B(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(G183gat), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT22), .B1(new_n215_), .B2(KEYINPUT78), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(KEYINPUT22), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n214_), .B(new_n216_), .C1(new_n217_), .C2(KEYINPUT78), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n215_), .A3(new_n214_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n222_), .A2(new_n223_), .B1(KEYINPUT24), .B2(new_n219_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n211_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n212_), .A2(KEYINPUT26), .ZN(new_n229_));
  OR2_X1    g028(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT30), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n209_), .B1(new_n234_), .B2(KEYINPUT80), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n235_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  OR2_X1    g040(.A1(new_n241_), .A2(KEYINPUT31), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT31), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n242_), .A2(KEYINPUT81), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n238_), .B(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G1gat), .B(G29gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252_));
  OR2_X1    g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G141gat), .ZN(new_n256_));
  INV_X1    g055(.A(G148gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n258_), .A2(KEYINPUT3), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT83), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n255_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n254_), .A2(KEYINPUT1), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(G155gat), .A3(G162gat), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n267_), .A2(new_n269_), .A3(new_n253_), .A4(KEYINPUT82), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(new_n268_), .A3(G155gat), .A4(G162gat), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n270_), .A2(new_n272_), .A3(new_n260_), .A4(new_n258_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n241_), .B1(new_n266_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n255_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n264_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n261_), .A2(new_n262_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n276_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n239_), .B(new_n240_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n273_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(KEYINPUT94), .A3(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n266_), .A2(new_n274_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT94), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n281_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n252_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(new_n275_), .B2(KEYINPUT4), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n251_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n283_), .A2(new_n286_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n288_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n295_), .B(new_n250_), .C1(new_n287_), .C2(new_n290_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n245_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299_));
  XOR2_X1   g098(.A(G8gat), .B(G36gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT91), .Z(new_n308_));
  OAI21_X1  g107(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n219_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT22), .B(G169gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n214_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n224_), .A2(new_n225_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT26), .B(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n227_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n211_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(G197gat), .B2(G204gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n323_), .B2(G197gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n323_), .B2(G197gat), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n324_), .B(new_n325_), .C1(new_n327_), .C2(KEYINPUT21), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT86), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n319_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n327_), .B(new_n330_), .C1(new_n329_), .C2(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n318_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT20), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n232_), .A2(new_n332_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n308_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT92), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n333_), .B(KEYINPUT20), .C1(new_n332_), .C2(new_n232_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(KEYINPUT92), .A3(new_n308_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n232_), .B2(new_n332_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n307_), .B1(new_n318_), .B2(new_n332_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n304_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n304_), .ZN(new_n349_));
  AOI211_X1 g148(.A(new_n349_), .B(new_n346_), .C1(new_n338_), .C2(new_n340_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n299_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n304_), .B(KEYINPUT99), .Z(new_n352_));
  NOR2_X1   g151(.A1(new_n339_), .A2(new_n308_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n318_), .A2(KEYINPUT98), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n328_), .A2(new_n331_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT98), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n313_), .B(new_n356_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n307_), .B1(new_n358_), .B2(new_n343_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n352_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n360_), .A2(KEYINPUT27), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n341_), .A2(new_n304_), .A3(new_n347_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n280_), .B2(new_n273_), .ZN(new_n366_));
  AND2_X1   g165(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(G228gat), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n369_), .A2(new_n370_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI22_X1  g172(.A1(new_n366_), .A2(new_n355_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n332_), .B(new_n372_), .C1(new_n284_), .C2(new_n365_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G78gat), .B(G106gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT88), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n374_), .A2(new_n375_), .A3(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n284_), .A2(new_n365_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G22gat), .B(G50gat), .Z(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT28), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n382_), .B(new_n384_), .ZN(new_n385_));
  AND4_X1   g184(.A1(KEYINPUT89), .A2(new_n380_), .A3(new_n381_), .A4(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n388_), .A2(new_n385_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n364_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n298_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n293_), .A2(new_n296_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n364_), .A2(new_n395_), .A3(KEYINPUT100), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT100), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n339_), .A2(KEYINPUT92), .A3(new_n308_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT92), .B1(new_n339_), .B2(new_n308_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n347_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n349_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n362_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n402_), .A2(new_n299_), .B1(new_n362_), .B2(new_n361_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n386_), .A2(new_n389_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(new_n297_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n397_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n396_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n296_), .A2(KEYINPUT33), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n294_), .A2(KEYINPUT4), .ZN(new_n409_));
  INV_X1    g208(.A(new_n290_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n295_), .A4(new_n250_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n283_), .A2(KEYINPUT96), .A3(new_n286_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT96), .B1(new_n283_), .B2(new_n286_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n289_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n288_), .B1(new_n275_), .B2(KEYINPUT4), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n417_), .B(new_n251_), .C1(new_n287_), .C2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n414_), .A2(new_n362_), .A3(new_n401_), .A4(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT97), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n348_), .A2(new_n350_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n414_), .A4(new_n419_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n400_), .B2(new_n425_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n394_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n421_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n404_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n407_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n393_), .B1(new_n432_), .B2(new_n245_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G229gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT72), .B(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G22gat), .ZN(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  INV_X1    g237(.A(G8gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G8gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n442_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G29gat), .B(G36gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G43gat), .B(G50gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n443_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n435_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n448_), .B(KEYINPUT15), .Z(new_n453_));
  OAI211_X1 g252(.A(new_n452_), .B(new_n434_), .C1(new_n445_), .C2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G113gat), .B(G141gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G169gat), .B(G197gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT101), .B1(new_n433_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n428_), .B1(new_n420_), .B2(KEYINPUT97), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n390_), .B1(new_n463_), .B2(new_n424_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT100), .B1(new_n364_), .B2(new_n395_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n403_), .A2(new_n397_), .A3(new_n405_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n245_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n392_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT101), .ZN(new_n470_));
  INV_X1    g269(.A(new_n461_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n462_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G85gat), .ZN(new_n474_));
  INV_X1    g273(.A(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT6), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n205_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n479_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n482_), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n480_), .A2(KEYINPUT6), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n488_), .B(new_n487_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n479_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n477_), .A2(KEYINPUT9), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n499_));
  OR2_X1    g298(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n486_), .A3(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n476_), .A2(KEYINPUT9), .A3(new_n477_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n448_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n505_), .A2(new_n506_), .B1(KEYINPUT35), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n508_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n488_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n481_), .A2(new_n483_), .ZN(new_n518_));
  AOI211_X1 g317(.A(KEYINPUT8), .B(new_n478_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n495_), .B1(new_n494_), .B2(new_n479_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n502_), .A2(new_n503_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT9), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(G85gat), .A3(G92gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n499_), .A2(KEYINPUT65), .A3(new_n502_), .A4(new_n503_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n521_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n527_), .A2(new_n528_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT66), .B1(new_n532_), .B2(new_n497_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n510_), .B(new_n514_), .C1(new_n534_), .C2(new_n453_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n530_), .B1(new_n521_), .B2(new_n529_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n497_), .A3(KEYINPUT66), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n453_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n513_), .B1(new_n538_), .B2(new_n509_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  OAI22_X1  g342(.A1(new_n540_), .A2(KEYINPUT71), .B1(KEYINPUT36), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n535_), .A2(new_n539_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(KEYINPUT36), .A3(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT37), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n552_), .A3(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n445_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n559_), .A3(KEYINPUT11), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  INV_X1    g360(.A(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G57gat), .ZN(new_n563_));
  INV_X1    g362(.A(G57gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(G64gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n565_), .A3(KEYINPUT11), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n558_), .A2(KEYINPUT11), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n560_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n557_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n557_), .A2(new_n569_), .ZN(new_n571_));
  XOR2_X1   g370(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT74), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G183gat), .B(G211gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT17), .ZN(new_n578_));
  AND4_X1   g377(.A1(new_n555_), .A2(new_n570_), .A3(new_n571_), .A4(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n570_), .A2(new_n571_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n555_), .B1(new_n580_), .B2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n570_), .A2(new_n571_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n504_), .B(new_n569_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(KEYINPUT67), .A3(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n569_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT12), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n505_), .A2(new_n595_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n594_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n589_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n588_), .B(KEYINPUT64), .ZN(new_n604_));
  INV_X1    g403(.A(new_n599_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT69), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  AND3_X1   g411(.A1(new_n602_), .A2(new_n606_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n602_), .B2(new_n606_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n587_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n612_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n588_), .A2(KEYINPUT67), .A3(new_n589_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT67), .B1(new_n588_), .B2(new_n589_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n596_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT12), .B1(new_n505_), .B2(new_n595_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT64), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n588_), .B(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n589_), .B1(new_n624_), .B2(new_n599_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n616_), .B1(new_n622_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n602_), .A2(new_n606_), .A3(new_n612_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT70), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n615_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT13), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n615_), .A2(new_n628_), .A3(KEYINPUT13), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n554_), .A2(new_n586_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n473_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n438_), .A3(new_n297_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n433_), .A2(new_n550_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n586_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n633_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n471_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT102), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n394_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n637_), .A2(new_n638_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n639_), .A2(new_n646_), .A3(new_n647_), .ZN(G1324gat));
  OAI21_X1  g447(.A(G8gat), .B1(new_n645_), .B2(new_n403_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n403_), .A2(G8gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n636_), .B2(new_n653_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n635_), .A2(KEYINPUT103), .A3(G8gat), .A4(new_n403_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n651_), .B(KEYINPUT40), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  OAI21_X1  g459(.A(G15gat), .B1(new_n645_), .B2(new_n245_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n635_), .A2(G15gat), .A3(new_n245_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n645_), .B2(new_n404_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n404_), .A2(G22gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n635_), .B2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n550_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n641_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n642_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n462_), .B2(new_n472_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n674_), .A2(G29gat), .A3(new_n394_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n641_), .A2(new_n461_), .A3(new_n633_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n469_), .B2(new_n554_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n554_), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT43), .B(new_n679_), .C1(new_n468_), .C2(new_n392_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT44), .B(new_n676_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n433_), .B2(new_n679_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n469_), .A2(new_n677_), .A3(new_n554_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(KEYINPUT106), .A3(KEYINPUT44), .A4(new_n676_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n676_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n394_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n691_), .A3(KEYINPUT107), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n688_), .B2(new_n691_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n675_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n403_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n688_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n672_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n403_), .A2(G36gat), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n433_), .A2(KEYINPUT101), .A3(new_n461_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n470_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n702_), .B(new_n703_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT45), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n673_), .A2(new_n708_), .A3(new_n703_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n696_), .A2(new_n697_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n698_), .B1(new_n701_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n698_), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n707_), .A2(new_n709_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n676_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n364_), .B1(new_n717_), .B2(KEYINPUT44), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n683_), .B2(new_n687_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n714_), .B(new_n715_), .C1(new_n719_), .C2(new_n699_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n713_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(new_n245_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n689_), .A2(new_n690_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n688_), .A2(G43gat), .A3(new_n722_), .A4(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT109), .B(G43gat), .Z(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(new_n674_), .B2(new_n245_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT47), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n724_), .A2(new_n727_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n673_), .B2(new_n390_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n688_), .A2(new_n723_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n390_), .A2(G50gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(G1331gat));
  NAND4_X1  g535(.A1(new_n640_), .A2(new_n461_), .A3(new_n633_), .A4(new_n641_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n394_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n469_), .A2(new_n461_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n554_), .A2(new_n586_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n633_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT110), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n740_), .A2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT112), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n297_), .A2(new_n564_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n738_), .B1(new_n745_), .B2(new_n746_), .ZN(G1332gat));
  OAI21_X1  g546(.A(G64gat), .B1(new_n737_), .B2(new_n403_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT48), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n364_), .A2(new_n562_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n745_), .B2(new_n750_), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n737_), .B2(new_n245_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT49), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n722_), .A2(new_n203_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n745_), .B2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n737_), .B2(new_n404_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n404_), .A2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n745_), .B2(new_n758_), .ZN(G1335gat));
  NAND3_X1  g558(.A1(new_n740_), .A2(new_n633_), .A3(new_n671_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n760_), .A2(G85gat), .A3(new_n394_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n641_), .A2(new_n642_), .A3(new_n471_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n686_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n474_), .B1(new_n763_), .B2(new_n297_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n761_), .A2(new_n764_), .ZN(G1336gat));
  NOR3_X1   g564(.A1(new_n760_), .A2(G92gat), .A3(new_n403_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n475_), .B1(new_n763_), .B2(new_n364_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n722_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n760_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n205_), .B1(new_n763_), .B2(new_n722_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n686_), .A2(new_n390_), .A3(new_n762_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n775_), .A2(new_n776_), .A3(G106gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n775_), .B2(G106gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n390_), .A2(new_n486_), .ZN(new_n779_));
  OAI22_X1  g578(.A1(new_n777_), .A2(new_n778_), .B1(new_n760_), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n782_));
  AND4_X1   g581(.A1(new_n782_), .A2(new_n741_), .A3(new_n642_), .A4(new_n461_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n634_), .B2(new_n461_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n461_), .A2(new_n613_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n602_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n594_), .A2(new_n598_), .A3(KEYINPUT55), .A4(new_n601_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n598_), .A2(new_n624_), .A3(new_n601_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n603_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n616_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n798_), .B(KEYINPUT56), .C1(new_n793_), .C2(new_n616_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n787_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n434_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n457_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n445_), .A2(new_n453_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n452_), .A2(new_n435_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n803_), .B(new_n804_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n458_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n613_), .A2(new_n614_), .A3(new_n587_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT70), .B1(new_n626_), .B2(new_n627_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n629_), .A2(KEYINPUT114), .A3(new_n809_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n670_), .B1(new_n802_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n808_), .A2(new_n613_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n616_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n794_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI221_X1 g623(.A(new_n820_), .B1(KEYINPUT115), .B2(KEYINPUT58), .C1(new_n794_), .C2(new_n821_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n554_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n550_), .A2(new_n818_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n813_), .B(new_n808_), .C1(new_n615_), .C2(new_n628_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT114), .B1(new_n629_), .B2(new_n809_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n821_), .B2(KEYINPUT113), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n786_), .B1(new_n834_), .B2(new_n800_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n827_), .B(new_n829_), .C1(new_n832_), .C2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT116), .B1(new_n837_), .B2(new_n828_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n819_), .B(new_n826_), .C1(new_n836_), .C2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n641_), .B1(new_n839_), .B2(KEYINPUT117), .ZN(new_n840_));
  INV_X1    g639(.A(new_n826_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n842_), .B(new_n843_), .C1(new_n838_), .C2(new_n836_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n785_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n245_), .A2(new_n394_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n391_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n839_), .A2(new_n586_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n785_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n848_), .A2(new_n471_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G113gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n836_), .A2(new_n838_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n550_), .B1(new_n832_), .B2(new_n835_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n826_), .B1(new_n857_), .B2(KEYINPUT57), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT117), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n586_), .A3(new_n844_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n850_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n847_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n461_), .A2(G113gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n855_), .B1(new_n863_), .B2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866_));
  INV_X1    g665(.A(G120gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n785_), .B1(new_n839_), .B2(new_n586_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n852_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n633_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n848_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n642_), .A2(KEYINPUT60), .ZN(new_n873_));
  MUX2_X1   g672(.A(KEYINPUT60), .B(new_n873_), .S(new_n867_), .Z(new_n874_));
  NAND3_X1  g673(.A1(new_n861_), .A2(new_n862_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n866_), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n870_), .B1(new_n863_), .B2(KEYINPUT59), .ZN(new_n878_));
  OAI211_X1 g677(.A(KEYINPUT118), .B(new_n875_), .C1(new_n878_), .C2(new_n867_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n848_), .A2(new_n641_), .A3(new_n853_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G127gat), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n586_), .A2(G127gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n863_), .B2(new_n883_), .ZN(G1342gat));
  NAND3_X1  g683(.A1(new_n848_), .A2(new_n554_), .A3(new_n853_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G134gat), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n670_), .A2(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n863_), .B2(new_n887_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n722_), .A2(new_n404_), .A3(new_n394_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n861_), .A2(new_n403_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n461_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n256_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n642_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n257_), .ZN(G1345gat));
  NOR2_X1   g693(.A1(new_n890_), .A2(new_n586_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT61), .B(G155gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n890_), .B2(new_n679_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n670_), .A2(G162gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n890_), .B2(new_n899_), .ZN(G1347gat));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n298_), .A2(new_n364_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n390_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n868_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n215_), .B1(new_n905_), .B2(new_n471_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n901_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(KEYINPUT119), .A3(new_n907_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n851_), .A2(new_n471_), .A3(new_n903_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G169gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(KEYINPUT120), .A3(KEYINPUT62), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n907_), .A3(G169gat), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n908_), .A2(new_n909_), .A3(new_n912_), .A4(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n851_), .A2(new_n917_), .A3(new_n903_), .ZN(new_n918_));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n868_), .B2(new_n904_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n471_), .A3(new_n311_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n916_), .A2(new_n921_), .ZN(G1348gat));
  NAND2_X1  g721(.A1(new_n861_), .A2(new_n404_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n923_), .A2(new_n214_), .A3(new_n642_), .A4(new_n902_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n642_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n925_));
  OR3_X1    g724(.A1(new_n925_), .A2(KEYINPUT122), .A3(G176gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(KEYINPUT122), .B1(new_n925_), .B2(G176gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n845_), .A2(new_n390_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n902_), .A2(new_n586_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G183gat), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  AOI211_X1 g730(.A(new_n227_), .B(new_n586_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT123), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n920_), .A2(new_n228_), .A3(new_n641_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n861_), .A2(new_n404_), .A3(new_n930_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n934_), .B(new_n935_), .C1(new_n936_), .C2(G183gat), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n937_), .ZN(G1350gat));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939_));
  INV_X1    g738(.A(G190gat), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(new_n920_), .B2(new_n554_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n550_), .A2(new_n315_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n939_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n943_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n679_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n945_), .B(KEYINPUT124), .C1(new_n940_), .C2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n944_), .A2(new_n947_), .ZN(G1351gat));
  NOR3_X1   g747(.A1(new_n722_), .A2(new_n403_), .A3(new_n395_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n861_), .A2(new_n471_), .A3(new_n949_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g750(.A(KEYINPUT125), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n861_), .A2(new_n949_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n642_), .ZN(new_n954_));
  INV_X1    g753(.A(G204gat), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n952_), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n954_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n957_));
  OAI211_X1 g756(.A(KEYINPUT125), .B(G204gat), .C1(new_n953_), .C2(new_n642_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n956_), .A2(new_n957_), .A3(new_n958_), .ZN(G1353gat));
  NAND2_X1  g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n641_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  XOR2_X1   g761(.A(new_n962_), .B(KEYINPUT126), .Z(new_n963_));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n953_), .A2(new_n961_), .A3(new_n965_), .ZN(new_n966_));
  OR2_X1    g765(.A1(new_n953_), .A2(new_n961_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n963_), .B(new_n964_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(G1354gat));
  OAI21_X1  g768(.A(G218gat), .B1(new_n953_), .B2(new_n679_), .ZN(new_n970_));
  OR2_X1    g769(.A1(new_n670_), .A2(G218gat), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n953_), .B2(new_n971_), .ZN(G1355gat));
endmodule


