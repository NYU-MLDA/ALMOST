//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n217_), .B2(new_n210_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n209_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  INV_X1    g021(.A(new_n208_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n207_), .A2(KEYINPUT65), .A3(new_n208_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n203_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT66), .A3(new_n219_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT66), .B1(new_n227_), .B2(new_n219_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n221_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT10), .B(G99gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n206_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n203_), .A4(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G29gat), .B(G36gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(G43gat), .B(G50gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n231_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n239_), .B(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT71), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n231_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT35), .ZN(new_n246_));
  INV_X1    g045(.A(new_n236_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n230_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT8), .A3(new_n228_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n249_), .B2(new_n221_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n245_), .B(new_n246_), .C1(new_n250_), .C2(new_n242_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G232gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n244_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT71), .B(new_n257_), .C1(new_n240_), .C2(new_n243_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G190gat), .B(G218gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT36), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n255_), .A2(new_n256_), .A3(new_n258_), .A4(new_n263_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n255_), .A2(new_n258_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n262_), .A2(KEYINPUT36), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT37), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n265_), .A2(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G57gat), .B(G64gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT11), .ZN(new_n280_));
  XOR2_X1   g079(.A(G71gat), .B(G78gat), .Z(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n280_), .A2(new_n281_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G231gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G1gat), .ZN(new_n287_));
  INV_X1    g086(.A(G8gat), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT14), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT74), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(KEYINPUT74), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G15gat), .B(G22gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT75), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n293_), .B(new_n295_), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n286_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT17), .ZN(new_n299_));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G183gat), .B(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  OR3_X1    g102(.A1(new_n298_), .A2(new_n299_), .A3(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(KEYINPUT17), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n277_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n231_), .A2(new_n236_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n284_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT12), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n284_), .ZN(new_n312_));
  INV_X1    g111(.A(G230gat), .ZN(new_n313_));
  INV_X1    g112(.A(G233gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT68), .B1(new_n312_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n318_));
  INV_X1    g117(.A(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n311_), .A2(new_n316_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(KEYINPUT67), .A3(new_n310_), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n309_), .A2(KEYINPUT67), .A3(new_n284_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n315_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G120gat), .B(G148gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(G176gat), .B(G204gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n321_), .A2(new_n324_), .A3(new_n330_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n332_), .A2(KEYINPUT13), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT13), .B1(new_n332_), .B2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n308_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT76), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G22gat), .B(G50gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G155gat), .B(G162gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT3), .ZN(new_n349_));
  INV_X1    g148(.A(G141gat), .ZN(new_n350_));
  INV_X1    g149(.A(G148gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n347_), .A2(new_n349_), .B1(new_n352_), .B2(KEYINPUT2), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT87), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n345_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n342_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(G155gat), .A3(G162gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT85), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT1), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT84), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n352_), .A2(new_n348_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n358_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n341_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n374_), .A3(new_n340_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT29), .B1(new_n358_), .B2(new_n370_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G197gat), .A2(G204gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G197gat), .A2(G204gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(KEYINPUT21), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT21), .ZN(new_n387_));
  INV_X1    g186(.A(new_n385_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n383_), .ZN(new_n389_));
  INV_X1    g188(.A(G218gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G211gat), .ZN(new_n391_));
  INV_X1    g190(.A(G211gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G218gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n386_), .B(new_n389_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n392_), .A2(G218gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n390_), .A2(G211gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT88), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n388_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n397_), .A2(new_n398_), .A3(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n395_), .A2(new_n396_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n386_), .A2(new_n389_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT89), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n382_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G228gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT90), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n382_), .A2(new_n411_), .A3(new_n408_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT91), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n416_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n415_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n414_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n381_), .A2(new_n418_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n415_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n380_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G1gat), .B(G29gat), .Z(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G57gat), .B(G85gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G127gat), .B(G134gat), .Z(new_n437_));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G127gat), .B(G134gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT83), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G113gat), .B(G120gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n358_), .B2(new_n370_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n436_), .B1(new_n446_), .B2(KEYINPUT4), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n368_), .A2(new_n369_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n443_), .A2(new_n444_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n345_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n356_), .B1(new_n345_), .B2(new_n353_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n448_), .B(new_n449_), .C1(new_n452_), .C2(new_n342_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n446_), .A2(new_n453_), .A3(KEYINPUT93), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT93), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n445_), .B(new_n455_), .C1(new_n358_), .C2(new_n370_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n447_), .B1(new_n457_), .B2(KEYINPUT4), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n436_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n434_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n435_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n461_), .B(new_n433_), .C1(new_n463_), .C2(new_n447_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT27), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G226gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n397_), .A2(new_n404_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G183gat), .A2(G190gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT78), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G183gat), .A3(G190gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n472_), .B1(new_n477_), .B2(KEYINPUT23), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(G183gat), .B2(G190gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n480_));
  INV_X1    g279(.A(G169gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT22), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G176gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT22), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT80), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G169gat), .A2(G176gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n486_), .B2(KEYINPUT80), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n479_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT25), .B(G183gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(G190gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(KEYINPUT24), .A3(new_n488_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n494_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n501_), .B1(G183gat), .B2(G190gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT23), .B1(new_n474_), .B2(new_n476_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n500_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n471_), .B1(new_n491_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G169gat), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n489_), .B1(new_n506_), .B2(new_n483_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n502_), .B1(new_n477_), .B2(new_n501_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(G183gat), .A2(G190gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n492_), .A2(new_n493_), .B1(new_n498_), .B2(new_n495_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n478_), .A2(new_n511_), .A3(new_n497_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT20), .B1(new_n513_), .B2(new_n408_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n470_), .B1(new_n505_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n491_), .A2(new_n504_), .A3(new_n471_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n408_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT20), .A4(new_n469_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G8gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT18), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G64gat), .B(G92gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n466_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n525_));
  AND4_X1   g324(.A1(KEYINPUT20), .A2(new_n516_), .A3(new_n470_), .A4(new_n517_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n513_), .B1(new_n409_), .B2(new_n405_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n505_), .ZN(new_n531_));
  OAI22_X1  g330(.A1(new_n503_), .A2(new_n502_), .B1(G183gat), .B2(G190gat), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n500_), .A2(new_n478_), .B1(new_n532_), .B2(new_n507_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n397_), .A2(new_n398_), .A3(new_n404_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n398_), .B1(new_n397_), .B2(new_n404_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n526_), .B1(new_n538_), .B2(new_n469_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n525_), .B1(new_n539_), .B2(new_n524_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n519_), .A2(new_n524_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n515_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n466_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n449_), .B(KEYINPUT31), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT82), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G71gat), .B(G99gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n491_), .A2(new_n504_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G227gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(G15gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT30), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n551_), .B(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT81), .B(G43gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n550_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n550_), .A2(new_n558_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n428_), .A2(new_n465_), .A3(new_n546_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n460_), .A2(new_n464_), .ZN(new_n563_));
  AOI211_X1 g362(.A(new_n563_), .B(new_n545_), .C1(new_n424_), .C2(new_n426_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n519_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n539_), .B2(new_n565_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT96), .B1(new_n465_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n464_), .B2(new_n460_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n464_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n457_), .A2(KEYINPUT4), .ZN(new_n574_));
  INV_X1    g373(.A(new_n446_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n436_), .B1(new_n575_), .B2(new_n462_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n433_), .B1(new_n457_), .B2(new_n436_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n543_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n447_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n581_), .A2(KEYINPUT33), .A3(new_n461_), .A4(new_n433_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n573_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n568_), .A2(new_n571_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n564_), .B1(new_n584_), .B2(new_n428_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n562_), .B1(new_n585_), .B2(new_n561_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n296_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n239_), .B(KEYINPUT77), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n296_), .A2(new_n242_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n589_), .A2(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G113gat), .B(G141gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n586_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n338_), .A2(KEYINPUT76), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n339_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n287_), .A3(new_n563_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT97), .Z(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT38), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(KEYINPUT38), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n274_), .B(KEYINPUT98), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n586_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n336_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n600_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n610_), .A2(new_n307_), .A3(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n465_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n606_), .A2(new_n607_), .A3(new_n615_), .ZN(G1324gat));
  AOI21_X1  g415(.A(new_n288_), .B1(new_n613_), .B2(new_n545_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT39), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n603_), .A2(new_n288_), .A3(new_n545_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g420(.A(new_n553_), .B1(new_n613_), .B2(new_n561_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n603_), .A2(new_n553_), .A3(new_n561_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n427_), .B(KEYINPUT99), .Z(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n613_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT42), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n603_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1327gat));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n586_), .A2(new_n633_), .A3(new_n277_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n583_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n636_));
  AOI211_X1 g435(.A(KEYINPUT96), .B(new_n567_), .C1(new_n464_), .C2(new_n460_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n428_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n427_), .A2(new_n546_), .A3(new_n465_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n561_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n562_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n635_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT100), .B(new_n562_), .C1(new_n585_), .C2(new_n561_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n272_), .A2(new_n276_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n642_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n648_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n648_), .B2(KEYINPUT43), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n634_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n307_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n610_), .A2(new_n652_), .A3(new_n611_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(KEYINPUT44), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n653_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n648_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n655_), .B1(new_n660_), .B2(new_n634_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n662_));
  OAI21_X1  g461(.A(new_n654_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(G29gat), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n465_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n610_), .A2(new_n652_), .A3(new_n274_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n601_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n563_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1328gat));
  OAI21_X1  g468(.A(G36gat), .B1(new_n663_), .B2(new_n546_), .ZN(new_n670_));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n671_), .A3(new_n545_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT104), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n674_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n670_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n670_), .A2(new_n675_), .A3(new_n676_), .A4(KEYINPUT46), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n561_), .ZN(new_n684_));
  INV_X1    g483(.A(G43gat), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n654_), .B(new_n686_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  INV_X1    g487(.A(new_n667_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n689_), .B2(new_n684_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n687_), .A2(new_n688_), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n688_), .B1(new_n687_), .B2(new_n690_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n687_), .A2(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT106), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n688_), .A3(new_n690_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n696_), .A3(new_n682_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1330gat));
  OAI21_X1  g497(.A(G50gat), .B1(new_n663_), .B2(new_n428_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n627_), .A2(G50gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT107), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n689_), .B2(new_n701_), .ZN(G1331gat));
  AND2_X1   g501(.A1(new_n586_), .A2(new_n611_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n308_), .A2(new_n610_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(KEYINPUT108), .B2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(KEYINPUT108), .B2(new_n704_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n563_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT109), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n336_), .A2(new_n307_), .A3(new_n600_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n609_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n465_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n708_), .A2(new_n712_), .ZN(G1332gat));
  OAI21_X1  g512(.A(G64gat), .B1(new_n710_), .B2(new_n546_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(G64gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n717_), .A3(new_n545_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1333gat));
  OAI21_X1  g518(.A(G71gat), .B1(new_n710_), .B2(new_n684_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT49), .ZN(new_n721_));
  INV_X1    g520(.A(G71gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(new_n722_), .A3(new_n561_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1334gat));
  OAI21_X1  g523(.A(G78gat), .B1(new_n710_), .B2(new_n627_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT111), .Z(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n627_), .A2(G78gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT112), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n706_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n727_), .A2(new_n728_), .A3(new_n731_), .ZN(G1335gat));
  NAND4_X1  g531(.A1(new_n703_), .A2(new_n610_), .A3(new_n307_), .A4(new_n271_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT113), .Z(new_n734_));
  AOI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n563_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT114), .Z(new_n736_));
  NAND3_X1  g535(.A1(new_n610_), .A2(new_n307_), .A3(new_n611_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n660_), .B2(new_n634_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n465_), .A2(new_n215_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(G1336gat));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n216_), .A3(new_n545_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n738_), .A2(new_n545_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n216_), .ZN(G1337gat));
  AOI21_X1  g542(.A(new_n205_), .B1(new_n738_), .B2(new_n561_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n561_), .A2(new_n232_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n734_), .B2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n206_), .A3(new_n427_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n738_), .A2(new_n427_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G106gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT52), .B(new_n206_), .C1(new_n738_), .C2(new_n427_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT53), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n748_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1339gat));
  INV_X1    g556(.A(G113gat), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n600_), .A2(new_n333_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n321_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n311_), .A2(KEYINPUT55), .A3(new_n320_), .A4(new_n316_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n310_), .A2(KEYINPUT12), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n310_), .A2(KEYINPUT12), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n312_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n315_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT115), .B(new_n312_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n762_), .B(new_n763_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n331_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n760_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n770_), .A2(new_n775_), .A3(new_n776_), .A4(new_n331_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n332_), .A2(new_n333_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n597_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n587_), .A2(new_n588_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n599_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n274_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n277_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n770_), .A2(new_n776_), .A3(new_n331_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n785_), .A2(new_n333_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n776_), .B1(new_n770_), .B2(new_n331_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT117), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n789_), .B1(new_n794_), .B2(KEYINPUT58), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT117), .B(new_n796_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n759_), .A2(new_n788_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n274_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n652_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n338_), .A2(new_n801_), .A3(new_n611_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT54), .B1(new_n337_), .B2(new_n600_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT118), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n795_), .A2(new_n797_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n774_), .A2(new_n777_), .B1(new_n779_), .B2(new_n785_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n759_), .B1(new_n807_), .B2(new_n271_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n799_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n307_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n802_), .A2(new_n803_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NOR4_X1   g613(.A1(new_n684_), .A2(new_n427_), .A3(new_n465_), .A4(new_n545_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n806_), .A2(KEYINPUT119), .A3(new_n808_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT119), .B1(new_n806_), .B2(new_n808_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n810_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n819_), .B2(new_n652_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n815_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n816_), .A2(KEYINPUT59), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n758_), .B1(new_n824_), .B2(new_n600_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n816_), .A2(G113gat), .A3(new_n611_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT120), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n820_), .A2(new_n823_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n600_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G113gat), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(new_n826_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n827_), .A2(new_n834_), .ZN(G1340gat));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n824_), .B2(new_n610_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(KEYINPUT60), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  AOI21_X1  g639(.A(G120gat), .B1(new_n610_), .B2(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n816_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n836_), .B1(new_n838_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n828_), .A2(new_n610_), .A3(new_n829_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G120gat), .ZN(new_n845_));
  INV_X1    g644(.A(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT121), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(G1341gat));
  INV_X1    g647(.A(new_n824_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G127gat), .B1(new_n849_), .B2(new_n307_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n307_), .A2(G127gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n816_), .B2(new_n851_), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n816_), .A2(new_n608_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(G134gat), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT122), .B(G134gat), .Z(new_n855_));
  NOR2_X1   g654(.A1(new_n789_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n824_), .B2(new_n856_), .ZN(G1343gat));
  NOR3_X1   g656(.A1(new_n428_), .A2(new_n465_), .A3(new_n545_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n805_), .A2(new_n814_), .A3(new_n684_), .A4(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n611_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n350_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n336_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n351_), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n859_), .A2(new_n307_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  NOR2_X1   g665(.A1(new_n859_), .A2(new_n608_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n647_), .A2(G162gat), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n867_), .A2(G162gat), .B1(new_n859_), .B2(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT123), .ZN(G1347gat));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n684_), .A2(new_n563_), .A3(new_n546_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n627_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n820_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n600_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n871_), .B1(new_n876_), .B2(G169gat), .ZN(new_n877_));
  AOI211_X1 g676(.A(KEYINPUT62), .B(new_n481_), .C1(new_n875_), .C2(new_n600_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n600_), .A2(new_n506_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT124), .Z(new_n880_));
  OAI22_X1  g679(.A1(new_n877_), .A2(new_n878_), .B1(new_n874_), .B2(new_n880_), .ZN(G1348gat));
  AOI21_X1  g680(.A(G176gat), .B1(new_n875_), .B2(new_n610_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n805_), .A2(new_n814_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n428_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT125), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n886_), .A3(new_n428_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n885_), .A2(new_n872_), .A3(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n336_), .A2(new_n483_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n882_), .B1(new_n888_), .B2(new_n889_), .ZN(G1349gat));
  NOR3_X1   g689(.A1(new_n874_), .A2(new_n307_), .A3(new_n492_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n885_), .A2(new_n652_), .A3(new_n872_), .A4(new_n887_), .ZN(new_n892_));
  INV_X1    g691(.A(G183gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1350gat));
  INV_X1    g693(.A(new_n493_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n608_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n875_), .A2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G190gat), .B1(new_n874_), .B2(new_n789_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT126), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n901_), .A3(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n428_), .A2(new_n563_), .A3(new_n546_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n805_), .A2(new_n814_), .A3(new_n684_), .A4(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n906_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G197gat), .B1(new_n909_), .B2(new_n600_), .ZN(new_n910_));
  INV_X1    g709(.A(G197gat), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n911_), .B(new_n611_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1352gat));
  INV_X1    g712(.A(new_n908_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n905_), .A2(new_n906_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n610_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G204gat), .ZN(new_n917_));
  INV_X1    g716(.A(G204gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n909_), .A2(new_n918_), .A3(new_n610_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1353gat));
  OR2_X1    g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n909_), .B2(new_n652_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT63), .B(G211gat), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n307_), .B(new_n923_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1354gat));
  NOR2_X1   g724(.A1(new_n608_), .A2(G218gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n909_), .A2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n789_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n390_), .B2(new_n928_), .ZN(G1355gat));
endmodule


