//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n205_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G229gat), .A2(G233gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n212_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n205_), .B2(new_n212_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n216_), .B1(new_n219_), .B2(new_n215_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G113gat), .B(G141gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G169gat), .B(G197gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n220_), .B(new_n225_), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT77), .ZN(new_n227_));
  AND3_X1   g026(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G183gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT78), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G183gat), .ZN(new_n234_));
  INV_X1    g033(.A(G190gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G169gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT26), .B(G190gat), .Z(new_n241_));
  NOR2_X1   g040(.A1(new_n233_), .A2(G183gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n231_), .A2(KEYINPUT78), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT25), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n241_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248_));
  INV_X1    g047(.A(G169gat), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT24), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n230_), .B(new_n251_), .C1(new_n252_), .C2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n240_), .B1(new_n247_), .B2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G71gat), .B(G99gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(G15gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G43gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n260_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266_));
  INV_X1    g065(.A(G120gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G113gat), .ZN(new_n268_));
  INV_X1    g067(.A(G113gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G120gat), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(new_n270_), .A3(KEYINPUT81), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT81), .B1(new_n268_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n266_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n269_), .A2(G120gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n267_), .A2(G113gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n266_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n268_), .A2(new_n270_), .A3(KEYINPUT81), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n273_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT82), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT31), .Z(new_n286_));
  AND2_X1   g085(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT83), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n265_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n265_), .A2(new_n289_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT21), .ZN(new_n293_));
  AND2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G197gat), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(KEYINPUT21), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n294_), .A2(new_n295_), .A3(new_n293_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308_));
  INV_X1    g107(.A(G141gat), .ZN(new_n309_));
  INV_X1    g108(.A(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G155gat), .B(G162gat), .Z(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G155gat), .ZN(new_n320_));
  INV_X1    g119(.A(G162gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT1), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G155gat), .A3(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n321_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G141gat), .B(G148gat), .Z(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(new_n328_), .ZN(new_n329_));
  AOI211_X1 g128(.A(KEYINPUT85), .B(new_n307_), .C1(KEYINPUT29), .C2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G78gat), .B(G106gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT86), .ZN(new_n332_));
  NAND2_X1  g131(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(G228gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n332_), .B(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n330_), .B(new_n337_), .Z(new_n338_));
  OR2_X1    g137(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT28), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G22gat), .B(G50gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n340_), .A2(new_n341_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n338_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n330_), .B(new_n337_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n342_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n252_), .B1(new_n254_), .B2(KEYINPUT89), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n253_), .A2(new_n351_), .A3(KEYINPUT24), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n251_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT26), .B(G190gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n353_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n230_), .B1(G183gat), .B2(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n239_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n303_), .A2(new_n306_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n360_), .B1(new_n373_), .B2(new_n245_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n254_), .A2(new_n252_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n358_), .A2(new_n375_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n374_), .A2(new_n376_), .B1(new_n239_), .B2(new_n237_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(new_n307_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n368_), .A2(new_n371_), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n256_), .B2(new_n367_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT88), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n363_), .A2(new_n365_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n384_), .B(KEYINPUT20), .C1(new_n256_), .C2(new_n367_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n379_), .B1(new_n386_), .B2(new_n371_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT91), .ZN(new_n389_));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n391_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(new_n383_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n374_), .A2(new_n376_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n307_), .A2(new_n398_), .A3(new_n240_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n384_), .B1(new_n399_), .B2(KEYINPUT20), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n397_), .A2(new_n371_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n371_), .B1(new_n368_), .B2(new_n378_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n396_), .B1(new_n404_), .B2(new_n395_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n408_), .A2(new_n410_), .ZN(new_n415_));
  OR3_X1    g214(.A1(new_n412_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n317_), .A2(new_n318_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n271_), .A2(new_n272_), .A3(new_n266_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(new_n283_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n285_), .A2(new_n329_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(KEYINPUT4), .A3(new_n423_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT92), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  AND4_X1   g231(.A1(new_n431_), .A2(new_n285_), .A3(new_n432_), .A4(new_n329_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n421_), .B2(new_n432_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n428_), .B(new_n430_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n435_), .B2(KEYINPUT93), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT92), .B1(new_n429_), .B2(KEYINPUT4), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n421_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n426_), .B1(new_n425_), .B2(KEYINPUT4), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n437_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n419_), .B1(new_n436_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n435_), .A2(KEYINPUT93), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n441_), .A3(new_n437_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n418_), .A4(new_n427_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n405_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n391_), .B(new_n392_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n371_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n377_), .B2(new_n307_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n382_), .B1(new_n451_), .B2(new_n384_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n449_), .B1(new_n452_), .B2(new_n381_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n448_), .B1(new_n453_), .B2(new_n379_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n371_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n379_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n394_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n426_), .B(new_n430_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n425_), .A2(new_n428_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n419_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n459_), .A2(new_n419_), .A3(KEYINPUT97), .A4(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n458_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n427_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n433_), .A2(new_n434_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n430_), .A2(new_n428_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n469_), .B2(new_n437_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(KEYINPUT33), .A3(new_n418_), .A4(new_n444_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n446_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n465_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT98), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n447_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n465_), .A2(new_n471_), .A3(KEYINPUT98), .A4(new_n473_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n349_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT99), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n457_), .A2(KEYINPUT27), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n452_), .A2(new_n449_), .A3(new_n381_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n394_), .B1(new_n481_), .B2(new_n402_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT27), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n453_), .A2(new_n448_), .A3(new_n379_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n394_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n484_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n448_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n457_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n349_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT100), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT100), .B1(new_n490_), .B2(new_n491_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n292_), .B1(new_n478_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n443_), .A2(new_n446_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n292_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n487_), .A2(new_n489_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n484_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT99), .B1(new_n501_), .B2(new_n488_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT101), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT101), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n483_), .A2(new_n504_), .A3(new_n487_), .A4(new_n489_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n349_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT102), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT102), .ZN(new_n509_));
  AOI211_X1 g308(.A(new_n509_), .B(new_n349_), .C1(new_n503_), .C2(new_n505_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n499_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n227_), .B1(new_n497_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G71gat), .B(G78gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT11), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n518_));
  INV_X1    g317(.A(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n517_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT64), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT10), .B(G99gat), .Z(new_n528_));
  INV_X1    g327(.A(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G85gat), .B(G92gat), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT9), .ZN(new_n532_));
  INV_X1    g331(.A(G85gat), .ZN(new_n533_));
  INV_X1    g332(.A(G92gat), .ZN(new_n534_));
  OR3_X1    g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT9), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n527_), .A2(new_n530_), .A3(new_n532_), .A4(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n531_), .B1(new_n539_), .B2(new_n526_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(KEYINPUT8), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n536_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n523_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n523_), .A2(new_n543_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n514_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT65), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT12), .B1(new_n523_), .B2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n523_), .A2(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n522_), .B(KEYINPUT67), .Z(new_n553_));
  OAI211_X1 g352(.A(KEYINPUT66), .B(new_n536_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .A4(KEYINPUT12), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n513_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT65), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n557_), .B(new_n514_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n547_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G120gat), .B(G148gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n547_), .A2(new_n556_), .A3(new_n558_), .A4(new_n564_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(KEYINPUT69), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT69), .B1(new_n566_), .B2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT13), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n567_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT69), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT13), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n568_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(new_n581_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT34), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n543_), .B2(new_n205_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n586_), .A2(new_n587_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n552_), .A2(new_n554_), .A3(new_n217_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT71), .ZN(new_n594_));
  INV_X1    g393(.A(new_n590_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n589_), .B(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n597_), .B2(new_n592_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n582_), .B(new_n583_), .C1(new_n594_), .C2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n593_), .B(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n592_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n590_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n601_), .A2(new_n603_), .A3(new_n581_), .A4(new_n580_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n599_), .A2(KEYINPUT37), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G127gat), .B(G155gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT17), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT74), .Z(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT72), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n212_), .B(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n553_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n553_), .A2(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT75), .ZN(new_n623_));
  INV_X1    g422(.A(new_n619_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(new_n523_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n523_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n614_), .A2(KEYINPUT17), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n625_), .A2(new_n615_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n577_), .A2(new_n609_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n512_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n207_), .A3(new_n498_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT38), .ZN(new_n634_));
  INV_X1    g433(.A(new_n226_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n577_), .A2(new_n635_), .A3(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n497_), .A2(new_n511_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT103), .B1(new_n638_), .B2(new_n605_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(KEYINPUT103), .A3(new_n605_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n498_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n634_), .A2(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n506_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n599_), .A2(new_n604_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n648_), .B(new_n649_), .C1(new_n497_), .C2(new_n511_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n647_), .B(new_n636_), .C1(new_n639_), .C2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G8gat), .B1(new_n651_), .B2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT39), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n642_), .A2(KEYINPUT104), .A3(new_n647_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n652_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(G8gat), .A4(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n632_), .A2(new_n208_), .A3(new_n647_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n660_), .A2(KEYINPUT40), .A3(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  OAI21_X1  g465(.A(G15gat), .B1(new_n643_), .B2(new_n292_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT41), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(KEYINPUT41), .ZN(new_n669_));
  INV_X1    g468(.A(new_n292_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n632_), .A2(new_n262_), .A3(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT105), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n669_), .A3(new_n672_), .ZN(G1326gat));
  OR3_X1    g472(.A1(new_n631_), .A2(G22gat), .A3(new_n507_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G22gat), .B1(new_n643_), .B2(new_n507_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT42), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT42), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679_));
  INV_X1    g478(.A(new_n577_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n649_), .A2(new_n629_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n512_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(G29gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n498_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n629_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n577_), .A2(new_n635_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n638_), .B2(new_n609_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n599_), .A2(KEYINPUT37), .A3(new_n604_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT37), .B1(new_n599_), .B2(new_n604_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n692_), .C1(new_n497_), .C2(new_n511_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n687_), .B(KEYINPUT44), .C1(new_n689_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n687_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n696_), .B2(KEYINPUT106), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n687_), .B(new_n698_), .C1(new_n689_), .C2(new_n693_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n695_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(new_n498_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n679_), .B(new_n685_), .C1(new_n701_), .C2(new_n684_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n684_), .B1(new_n700_), .B2(new_n498_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n685_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT107), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n506_), .A2(G36gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n683_), .B2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n683_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n709_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n696_), .A2(KEYINPUT106), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n699_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n647_), .A3(new_n694_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n711_), .A2(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT46), .B(new_n713_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  AOI21_X1  g522(.A(G43gat), .B1(new_n683_), .B2(new_n670_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n670_), .A2(G43gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n700_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n683_), .B2(new_n349_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n349_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n700_), .B2(new_n730_), .ZN(G1331gat));
  AOI211_X1 g530(.A(new_n226_), .B(new_n680_), .C1(new_n497_), .C2(new_n511_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n690_), .A2(new_n691_), .A3(new_n629_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G57gat), .B1(new_n734_), .B2(new_n498_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n639_), .A2(new_n650_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n577_), .A2(new_n686_), .A3(new_n227_), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n736_), .A2(KEYINPUT110), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT110), .B1(new_n736_), .B2(new_n737_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT111), .B(G57gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n644_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(KEYINPUT112), .A3(new_n742_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n735_), .B1(new_n745_), .B2(new_n746_), .ZN(G1332gat));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n734_), .A2(new_n748_), .A3(new_n647_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n738_), .A2(new_n647_), .A3(new_n739_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G64gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G64gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n734_), .A2(new_n755_), .A3(new_n670_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n738_), .A2(new_n670_), .A3(new_n739_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G71gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1334gat));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n734_), .A2(new_n762_), .A3(new_n349_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n738_), .A2(new_n349_), .A3(new_n739_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G78gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G78gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1335gat));
  NOR3_X1   g567(.A1(new_n680_), .A2(new_n226_), .A3(new_n686_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n644_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n732_), .A2(new_n772_), .A3(new_n682_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n732_), .B2(new_n682_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n498_), .A2(new_n533_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n771_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT114), .ZN(G1336gat));
  OAI21_X1  g577(.A(G92gat), .B1(new_n770_), .B2(new_n506_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n647_), .A2(new_n534_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n775_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT115), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n770_), .B2(new_n292_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n670_), .A2(new_n528_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n775_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g585(.A(G106gat), .B1(new_n770_), .B2(new_n507_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n788_));
  AND2_X1   g587(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n788_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n529_), .B(new_n349_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n790_), .A2(new_n795_), .A3(new_n791_), .A4(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n508_), .A2(new_n510_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n292_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n513_), .B1(new_n550_), .B2(new_n555_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n556_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n550_), .A2(new_n555_), .A3(KEYINPUT55), .A4(new_n513_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n565_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT56), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n220_), .A2(new_n223_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n213_), .A2(new_n215_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n219_), .B(KEYINPUT117), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n214_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n807_), .B1(new_n810_), .B2(new_n223_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n812_), .A3(new_n565_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n806_), .A2(new_n567_), .A3(new_n811_), .A4(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(KEYINPUT58), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT118), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n609_), .B1(new_n815_), .B2(KEYINPUT58), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n806_), .A2(new_n226_), .A3(new_n567_), .A4(new_n813_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n574_), .A2(new_n568_), .A3(new_n811_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT57), .B1(new_n826_), .B2(new_n605_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n649_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n686_), .B1(new_n823_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n733_), .A2(new_n571_), .A3(new_n576_), .A4(new_n227_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n799_), .B(new_n498_), .C1(new_n831_), .C2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n226_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n827_), .A2(new_n829_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n821_), .B1(new_n819_), .B2(new_n817_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n629_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n832_), .B(KEYINPUT54), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n644_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(KEYINPUT59), .A3(new_n799_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n835_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT119), .B(G113gat), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n227_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n837_), .B1(new_n846_), .B2(new_n848_), .ZN(G1340gat));
  XOR2_X1   g648(.A(KEYINPUT120), .B(G120gat), .Z(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n680_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n836_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n850_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n680_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n850_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n852_), .B(KEYINPUT121), .C1(new_n853_), .C2(new_n850_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1341gat));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n836_), .A2(new_n859_), .A3(new_n686_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n629_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g661(.A(G134gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n836_), .A2(new_n863_), .A3(new_n649_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n692_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n292_), .A2(new_n349_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n647_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n498_), .B(new_n868_), .C1(new_n831_), .C2(new_n834_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n635_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n309_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n680_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n310_), .ZN(G1345gat));
  OAI21_X1  g672(.A(KEYINPUT122), .B1(new_n869_), .B2(new_n629_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n842_), .A2(new_n875_), .A3(new_n686_), .A4(new_n868_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n878_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n874_), .A2(new_n876_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n880_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n869_), .B2(new_n692_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n649_), .A2(new_n321_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n869_), .B2(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT124), .ZN(G1347gat));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n840_), .A2(new_n841_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n893_), .A2(new_n647_), .A3(new_n507_), .A4(new_n499_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n635_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT22), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n892_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G169gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n249_), .B1(new_n895_), .B2(new_n892_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(new_n899_), .ZN(G1348gat));
  NOR2_X1   g699(.A1(new_n894_), .A2(new_n680_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n250_), .ZN(G1349gat));
  NAND2_X1  g701(.A1(new_n232_), .A2(new_n234_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n894_), .A2(new_n629_), .ZN(new_n904_));
  MUX2_X1   g703(.A(new_n903_), .B(new_n361_), .S(new_n904_), .Z(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n894_), .B2(new_n692_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n649_), .A2(new_n360_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n894_), .B2(new_n907_), .ZN(G1351gat));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n867_), .A2(new_n498_), .A3(new_n506_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n893_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n226_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n909_), .B1(new_n913_), .B2(new_n297_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n297_), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n912_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n226_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(G1352gat));
  NOR2_X1   g716(.A1(new_n911_), .A2(new_n680_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n298_), .ZN(G1353gat));
  AOI21_X1  g718(.A(new_n629_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n912_), .A2(new_n920_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n923_));
  OAI22_X1  g722(.A1(new_n922_), .A2(new_n923_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n924_), .A2(new_n928_), .ZN(G1354gat));
  AND3_X1   g728(.A1(new_n912_), .A2(G218gat), .A3(new_n609_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n911_), .A2(KEYINPUT127), .A3(new_n605_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(G218gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT127), .B1(new_n911_), .B2(new_n605_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n930_), .B1(new_n932_), .B2(new_n933_), .ZN(G1355gat));
endmodule


