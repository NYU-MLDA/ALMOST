//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n971_,
    new_n972_, new_n974_, new_n975_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n998_, new_n999_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G43gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT80), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT81), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G71gat), .B(G99gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n208_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT23), .ZN(new_n214_));
  OR2_X1    g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT26), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT79), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n223_), .B(new_n224_), .C1(new_n228_), .C2(KEYINPUT79), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n217_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n220_), .A2(new_n229_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n212_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT31), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n205_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(new_n241_), .A3(new_n204_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OR3_X1    g046(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT86), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .A4(KEYINPUT84), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261_));
  OAI22_X1  g060(.A1(new_n261_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n255_), .A2(new_n256_), .A3(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n254_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n253_), .A2(KEYINPUT85), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT86), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n252_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n258_), .A2(new_n259_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n267_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n250_), .A2(KEYINPUT1), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n250_), .A2(KEYINPUT1), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n280_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n276_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n274_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n205_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n256_), .B1(new_n255_), .B2(new_n264_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n266_), .A2(KEYINPUT86), .A3(new_n272_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n288_), .B2(new_n252_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n204_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(KEYINPUT4), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G225gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n284_), .A2(new_n294_), .A3(new_n205_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n285_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G29gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT0), .ZN(new_n300_));
  INV_X1    g099(.A(G57gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G85gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n297_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n247_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n289_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT28), .ZN(new_n313_));
  XOR2_X1   g112(.A(G22gat), .B(G50gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  OR2_X1    g118(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  NAND2_X1  g120(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(G197gat), .A4(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n325_));
  INV_X1    g124(.A(G197gat), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT88), .B1(new_n326_), .B2(G204gat), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n319_), .B(new_n323_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G211gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(G218gat), .ZN(new_n331_));
  INV_X1    g130(.A(G218gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(G211gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT89), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(G211gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(G218gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(G197gat), .B1(new_n320_), .B2(new_n322_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n326_), .A2(G204gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT21), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n329_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT90), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n326_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n341_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n348_), .A2(KEYINPUT21), .B1(new_n334_), .B2(new_n338_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT90), .A3(new_n329_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n339_), .A2(new_n319_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n323_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n284_), .B2(KEYINPUT29), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n251_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(KEYINPUT29), .C1(new_n358_), .C2(new_n282_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n355_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n362_));
  INV_X1    g161(.A(G228gat), .ZN(new_n363_));
  INV_X1    g162(.A(G233gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n345_), .A2(new_n350_), .B1(new_n353_), .B2(new_n352_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT91), .B1(new_n289_), .B2(new_n311_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n359_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT92), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n355_), .A3(new_n370_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n318_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n374_), .ZN(new_n376_));
  AOI211_X1 g175(.A(new_n376_), .B(new_n317_), .C1(new_n366_), .C2(new_n371_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n316_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n362_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n369_), .A2(KEYINPUT92), .A3(new_n370_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n317_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n374_), .A3(new_n318_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n315_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n222_), .A2(new_n226_), .A3(KEYINPUT95), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT95), .B1(new_n222_), .B2(new_n226_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n224_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT96), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n220_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n224_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n391_), .A2(new_n398_), .A3(new_n393_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT96), .B1(new_n399_), .B2(new_n219_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n233_), .A2(KEYINPUT97), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n233_), .A2(KEYINPUT97), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n235_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n390_), .B1(new_n355_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n367_), .B2(new_n236_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AND4_X1   g207(.A1(KEYINPUT90), .A2(new_n329_), .A3(new_n339_), .A4(new_n342_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT90), .B1(new_n349_), .B2(new_n329_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n236_), .B(new_n354_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT20), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT94), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT94), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n414_), .A3(KEYINPUT20), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n351_), .A2(new_n354_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n418_), .B2(new_n389_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT18), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n412_), .A2(KEYINPUT94), .B1(new_n355_), .B2(new_n405_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n390_), .A3(new_n415_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n367_), .B(new_n404_), .C1(new_n219_), .C2(new_n399_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n389_), .B1(new_n428_), .B2(new_n407_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n424_), .B(KEYINPUT27), .C1(new_n430_), .C2(new_n423_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n390_), .B1(new_n425_), .B2(new_n415_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  INV_X1    g232(.A(new_n423_), .ZN(new_n434_));
  NOR4_X1   g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n408_), .A4(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT98), .B1(new_n419_), .B2(new_n423_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n424_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n437_), .B2(KEYINPUT27), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n310_), .A2(new_n386_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT102), .ZN(new_n440_));
  INV_X1    g239(.A(new_n308_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n378_), .A2(new_n384_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n378_), .A2(new_n384_), .A3(new_n441_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n432_), .A2(new_n408_), .A3(new_n434_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n423_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT27), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n419_), .A2(KEYINPUT98), .A3(new_n423_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n408_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n411_), .A2(new_n414_), .A3(KEYINPUT20), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n414_), .B1(new_n411_), .B2(KEYINPUT20), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n416_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n450_), .B1(new_n453_), .B2(new_n390_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n433_), .B1(new_n454_), .B2(new_n434_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n449_), .B1(new_n455_), .B2(new_n445_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n448_), .B1(new_n456_), .B2(new_n447_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n444_), .A2(new_n457_), .A3(KEYINPUT102), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n307_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n295_), .A2(new_n292_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n306_), .B1(new_n461_), .B2(new_n291_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n285_), .A2(KEYINPUT99), .A3(new_n290_), .ZN(new_n463_));
  AOI21_X1  g262(.A(KEYINPUT99), .B1(new_n285_), .B2(new_n290_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n293_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n307_), .A2(new_n459_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n460_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n436_), .A2(new_n424_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n449_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n423_), .A2(KEYINPUT32), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT101), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n472_), .A2(new_n473_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT101), .B1(new_n430_), .B2(new_n471_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT100), .B1(new_n419_), .B2(new_n471_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n419_), .A2(KEYINPUT100), .A3(new_n471_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n474_), .B(new_n475_), .C1(new_n476_), .C2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n470_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n385_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n443_), .A2(new_n458_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n439_), .B1(new_n481_), .B2(new_n247_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G71gat), .B(G78gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(KEYINPUT11), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT69), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G57gat), .B(G64gat), .Z(new_n488_));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(KEYINPUT69), .A3(new_n483_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n489_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n487_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n487_), .B2(new_n491_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G85gat), .B(G92gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT68), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  OAI22_X1  g302(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n502_), .B(new_n503_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n499_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n510_), .B(new_n499_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT66), .B(KEYINPUT9), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(new_n517_), .B2(new_n497_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(G85gat), .A4(G92gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n512_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n496_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G230gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT73), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n496_), .A2(new_n525_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT12), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n494_), .A2(new_n495_), .A3(new_n532_), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n517_), .A2(new_n497_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n522_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .A4(new_n516_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT72), .B1(new_n518_), .B2(new_n522_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n512_), .A2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n531_), .A2(new_n532_), .B1(new_n533_), .B2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n485_), .A2(new_n486_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT69), .B1(new_n490_), .B2(new_n483_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n492_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n487_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n523_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n529_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT73), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n530_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT70), .B1(new_n496_), .B2(new_n525_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n553_), .A3(new_n547_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n531_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(KEYINPUT71), .A3(new_n529_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT71), .B1(new_n555_), .B2(new_n529_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  NOR3_X1   g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT13), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT13), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n568_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G1gat), .B(G8gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT76), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n572_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G29gat), .B(G36gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G43gat), .B(G50gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G43gat), .B(G50gat), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n579_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n578_), .B(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n578_), .A2(new_n585_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n585_), .B(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n593_), .B2(new_n578_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT78), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n590_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n570_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n482_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n593_), .B1(new_n512_), .B2(new_n539_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  OAI22_X1  g411(.A1(new_n525_), .A2(new_n586_), .B1(KEYINPUT35), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n612_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n610_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n619_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT75), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n623_), .B(new_n627_), .C1(new_n619_), .C2(new_n624_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n625_), .A2(new_n626_), .A3(KEYINPUT37), .A4(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n578_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(new_n546_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G127gat), .B(G155gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT16), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT77), .B1(new_n640_), .B2(KEYINPUT17), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n640_), .A2(KEYINPUT17), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n633_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n609_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n574_), .A3(new_n308_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n481_), .A2(new_n247_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n439_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n625_), .A2(new_n628_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(KEYINPUT104), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657_));
  INV_X1    g456(.A(new_n655_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n482_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n607_), .A2(new_n645_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n661_), .A2(new_n441_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n651_), .B1(new_n574_), .B2(new_n663_), .ZN(G1324gat));
  XOR2_X1   g463(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n665_));
  NOR2_X1   g464(.A1(new_n662_), .A2(new_n457_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT106), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n575_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT104), .B1(new_n654_), .B2(new_n655_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n482_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT106), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(KEYINPUT39), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n457_), .A2(G8gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n648_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n648_), .A2(KEYINPUT105), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT39), .B1(new_n670_), .B2(new_n674_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n665_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n670_), .A2(new_n674_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n665_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n687_), .A2(new_n675_), .A3(new_n681_), .A4(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n684_), .A2(new_n689_), .ZN(G1325gat));
  INV_X1    g489(.A(new_n247_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n660_), .A2(new_n607_), .A3(new_n645_), .A4(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G15gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT41), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n692_), .A2(new_n695_), .A3(G15gat), .ZN(new_n696_));
  INV_X1    g495(.A(G15gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n648_), .A2(new_n697_), .A3(new_n691_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n694_), .A2(KEYINPUT108), .A3(new_n696_), .A4(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1326gat));
  INV_X1    g502(.A(G22gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n648_), .A2(new_n704_), .A3(new_n386_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n661_), .A2(new_n662_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n386_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n708_), .B2(G22gat), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT42), .B(new_n704_), .C1(new_n707_), .C2(new_n386_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(G1327gat));
  NOR2_X1   g510(.A1(new_n655_), .A2(new_n645_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n609_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n714_), .B2(new_n308_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n470_), .A2(new_n478_), .B1(new_n384_), .B2(new_n378_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n438_), .A2(new_n442_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(KEYINPUT102), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n691_), .B1(new_n719_), .B2(new_n443_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n716_), .B(new_n633_), .C1(new_n720_), .C2(new_n439_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n633_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n482_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n724_), .A2(KEYINPUT44), .A3(new_n607_), .A4(new_n646_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(G29gat), .A3(new_n308_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n646_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n608_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n715_), .B1(new_n726_), .B2(new_n729_), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n608_), .B(new_n645_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n457_), .B1(new_n733_), .B2(KEYINPUT44), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n734_), .B2(new_n729_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n714_), .A2(new_n732_), .A3(new_n438_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n731_), .B1(new_n735_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n733_), .A2(KEYINPUT44), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n725_), .A2(new_n438_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G36gat), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n736_), .B(KEYINPUT45), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n743_), .A3(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n744_), .ZN(G1329gat));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(G43gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n713_), .B2(new_n247_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n725_), .A2(G43gat), .A3(new_n691_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n740_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT47), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n747_), .C1(new_n748_), .C2(new_n740_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1330gat));
  AOI21_X1  g552(.A(G50gat), .B1(new_n714_), .B2(new_n386_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n725_), .A2(G50gat), .A3(new_n386_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n729_), .ZN(G1331gat));
  OR2_X1    g555(.A1(new_n567_), .A2(new_n569_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n605_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n482_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(new_n647_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n301_), .A3(new_n308_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n645_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n308_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n765_), .B2(new_n301_), .ZN(G1332gat));
  INV_X1    g565(.A(G64gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n761_), .A2(new_n767_), .A3(new_n438_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n764_), .B2(new_n438_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n769_), .A2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n761_), .A2(new_n774_), .A3(new_n691_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n764_), .A2(new_n691_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G71gat), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT49), .B(new_n774_), .C1(new_n764_), .C2(new_n691_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT110), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n775_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1334gat));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n761_), .A2(new_n785_), .A3(new_n386_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n764_), .B2(new_n386_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n788_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1335gat));
  AND2_X1   g590(.A1(new_n760_), .A2(new_n712_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G85gat), .B1(new_n792_), .B2(new_n308_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT111), .Z(new_n794_));
  NOR2_X1   g593(.A1(new_n728_), .A2(new_n759_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n441_), .A2(new_n303_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(G1336gat));
  INV_X1    g596(.A(G92gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n792_), .A2(new_n798_), .A3(new_n438_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n728_), .A2(new_n457_), .A3(new_n759_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n798_), .ZN(G1337gat));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n724_), .A2(new_n646_), .A3(new_n691_), .A4(new_n758_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G99gat), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n691_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n792_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n807_), .B2(KEYINPUT51), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n803_), .A2(G99gat), .B1(new_n792_), .B2(new_n805_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(KEYINPUT113), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT112), .B1(new_n807_), .B2(KEYINPUT51), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n809_), .A2(new_n813_), .A3(new_n810_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n808_), .B(new_n811_), .C1(new_n812_), .C2(new_n814_), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n792_), .A2(new_n514_), .A3(new_n386_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n724_), .A2(new_n646_), .A3(new_n386_), .A4(new_n758_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(G106gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n817_), .B2(G106gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT53), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(new_n816_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1339gat));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n594_), .A2(KEYINPUT117), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n594_), .A2(KEYINPUT117), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n588_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n599_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n601_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n562_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n532_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n496_), .A2(new_n540_), .A3(KEYINPUT12), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n552_), .A2(new_n835_), .A3(new_n836_), .A4(new_n554_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n529_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT116), .A3(new_n529_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n835_), .B(new_n836_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n548_), .A2(new_n549_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n840_), .A2(new_n841_), .B1(KEYINPUT55), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT115), .B(new_n846_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n834_), .B1(new_n845_), .B2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(KEYINPUT56), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n854_), .B(new_n834_), .C1(new_n845_), .C2(new_n851_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n564_), .B(new_n833_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n722_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n856_), .B2(new_n857_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n850_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n551_), .B2(new_n846_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n841_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT116), .B1(new_n837_), .B2(new_n529_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n864_), .A2(new_n865_), .B1(new_n846_), .B2(new_n551_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n562_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n854_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n852_), .A2(KEYINPUT56), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n563_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(KEYINPUT58), .A4(new_n833_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n859_), .B1(new_n860_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n833_), .A2(new_n566_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n870_), .B2(new_n605_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n874_), .B1(new_n877_), .B2(new_n658_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n564_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n879_), .B2(new_n606_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT57), .A3(new_n655_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n646_), .B1(new_n873_), .B2(new_n882_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n633_), .A2(new_n605_), .A3(new_n646_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n757_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT114), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n757_), .A2(new_n884_), .A3(new_n888_), .A4(new_n885_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n884_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n890_), .B2(new_n570_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n887_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n883_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n457_), .A2(new_n308_), .A3(new_n691_), .A4(new_n385_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT120), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n826_), .B1(new_n897_), .B2(new_n606_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n898_), .A2(KEYINPUT121), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n605_), .A2(G113gat), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n894_), .A2(new_n896_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(KEYINPUT59), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n897_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n900_), .B1(new_n902_), .B2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n898_), .A2(KEYINPUT121), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n899_), .A2(new_n905_), .A3(new_n906_), .ZN(G1340gat));
  XNOR2_X1  g706(.A(new_n897_), .B(KEYINPUT59), .ZN(new_n908_));
  OAI21_X1  g707(.A(G120gat), .B1(new_n908_), .B2(new_n757_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n910_));
  INV_X1    g709(.A(G120gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n570_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n901_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n901_), .A2(KEYINPUT122), .A3(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n909_), .A2(new_n918_), .ZN(G1341gat));
  OAI21_X1  g718(.A(G127gat), .B1(new_n908_), .B2(new_n646_), .ZN(new_n920_));
  OR3_X1    g719(.A1(new_n897_), .A2(G127gat), .A3(new_n646_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1342gat));
  OAI21_X1  g721(.A(G134gat), .B1(new_n908_), .B2(new_n722_), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n897_), .A2(G134gat), .A3(new_n655_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1343gat));
  NAND2_X1  g724(.A1(new_n860_), .A2(new_n872_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n858_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(new_n878_), .A3(new_n881_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n892_), .B1(new_n928_), .B2(new_n646_), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n438_), .A2(new_n691_), .A3(new_n385_), .A4(new_n441_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT123), .B1(new_n929_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n878_), .A2(new_n881_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n645_), .B1(new_n934_), .B2(new_n927_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n933_), .B(new_n930_), .C1(new_n935_), .C2(new_n892_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n932_), .A2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n605_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n570_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g740(.A1(new_n937_), .A2(new_n645_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT61), .B(G155gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1346gat));
  AOI21_X1  g743(.A(new_n933_), .B1(new_n894_), .B2(new_n930_), .ZN(new_n945_));
  AOI211_X1 g744(.A(KEYINPUT123), .B(new_n931_), .C1(new_n883_), .C2(new_n893_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n658_), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948_));
  INV_X1    g747(.A(G162gat), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n655_), .B1(new_n932_), .B2(new_n936_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT124), .B1(new_n951_), .B2(G162gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n937_), .A2(G162gat), .A3(new_n633_), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n950_), .A2(new_n952_), .A3(new_n953_), .ZN(G1347gat));
  NOR3_X1   g753(.A1(new_n310_), .A2(new_n386_), .A3(new_n457_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n894_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n894_), .A2(new_n955_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(KEYINPUT125), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n958_), .A2(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n961_), .A2(new_n605_), .A3(new_n230_), .ZN(new_n962_));
  OAI21_X1  g761(.A(G169gat), .B1(new_n959_), .B2(new_n606_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n963_), .A2(KEYINPUT62), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(KEYINPUT62), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n962_), .B1(new_n964_), .B2(new_n965_), .ZN(G1348gat));
  OAI21_X1  g765(.A(G176gat), .B1(new_n959_), .B2(new_n757_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n961_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n570_), .A2(new_n231_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n967_), .B1(new_n968_), .B2(new_n969_), .ZN(G1349gat));
  AOI21_X1  g769(.A(G183gat), .B1(new_n956_), .B2(new_n645_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n646_), .A2(new_n224_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(new_n961_), .B2(new_n972_), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n658_), .A2(new_n394_), .A3(new_n392_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n722_), .B1(new_n958_), .B2(new_n960_), .ZN(new_n975_));
  OAI22_X1  g774(.A1(new_n968_), .A2(new_n974_), .B1(new_n975_), .B2(new_n221_), .ZN(G1351gat));
  NOR3_X1   g775(.A1(new_n457_), .A2(new_n442_), .A3(new_n691_), .ZN(new_n977_));
  AND2_X1   g776(.A1(new_n894_), .A2(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(new_n605_), .ZN(new_n979_));
  AND3_X1   g778(.A1(new_n979_), .A2(KEYINPUT126), .A3(new_n326_), .ZN(new_n980_));
  AOI21_X1  g779(.A(KEYINPUT126), .B1(new_n979_), .B2(new_n326_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n979_), .A2(new_n326_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n980_), .A2(new_n981_), .A3(new_n982_), .ZN(G1352gat));
  NAND2_X1  g782(.A1(new_n894_), .A2(new_n977_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(new_n757_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n985_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n986_));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n987_));
  INV_X1    g786(.A(G204gat), .ZN(new_n988_));
  OAI211_X1 g787(.A(new_n986_), .B(new_n987_), .C1(new_n988_), .C2(new_n985_), .ZN(new_n989_));
  NOR4_X1   g788(.A1(new_n984_), .A2(new_n757_), .A3(new_n325_), .A4(new_n324_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n988_), .B1(new_n978_), .B2(new_n570_), .ZN(new_n991_));
  OAI21_X1  g790(.A(KEYINPUT127), .B1(new_n990_), .B2(new_n991_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n989_), .A2(new_n992_), .ZN(G1353gat));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n994_));
  OAI211_X1 g793(.A(new_n978_), .B(new_n645_), .C1(new_n994_), .C2(new_n330_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n994_), .A2(new_n330_), .ZN(new_n996_));
  XNOR2_X1  g795(.A(new_n995_), .B(new_n996_), .ZN(G1354gat));
  NAND3_X1  g796(.A1(new_n978_), .A2(new_n332_), .A3(new_n658_), .ZN(new_n998_));
  OAI21_X1  g797(.A(G218gat), .B1(new_n984_), .B2(new_n722_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n998_), .A2(new_n999_), .ZN(G1355gat));
endmodule


