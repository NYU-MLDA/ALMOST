//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n572_, new_n573_, new_n574_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n208_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT75), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n212_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n208_), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n217_), .B(KEYINPUT76), .Z(new_n222_));
  AND3_X1   g021(.A1(new_n221_), .A2(new_n213_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G113gat), .B(G141gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G169gat), .B(G197gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n228_), .B(new_n229_), .Z(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n219_), .A2(new_n225_), .A3(new_n226_), .A4(new_n230_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n242_));
  INV_X1    g041(.A(G183gat), .ZN(new_n243_));
  INV_X1    g042(.A(G190gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT81), .ZN(new_n246_));
  NOR2_X1   g045(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G169gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G169gat), .ZN(new_n250_));
  INV_X1    g049(.A(G176gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(KEYINPUT24), .A3(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n255_), .B1(new_n239_), .B2(new_n237_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n243_), .A2(KEYINPUT25), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n244_), .A2(KEYINPUT26), .ZN(new_n259_));
  AOI22_X1  g058(.A1(KEYINPUT78), .A2(new_n258_), .B1(new_n259_), .B2(KEYINPUT79), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(KEYINPUT79), .B2(new_n259_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n243_), .A2(KEYINPUT25), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n244_), .A2(KEYINPUT26), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n262_), .B(new_n263_), .C1(new_n258_), .C2(KEYINPUT78), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n254_), .B(new_n256_), .C1(new_n261_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n249_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT21), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT21), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n266_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G226gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT25), .B(G183gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n254_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT86), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n242_), .A2(new_n255_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT87), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(KEYINPUT87), .A3(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n237_), .A2(new_n239_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT88), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n274_), .B1(new_n248_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n275_), .A2(KEYINPUT20), .A3(new_n278_), .A4(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G8gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT18), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G64gat), .B(G92gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT32), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT20), .B1(new_n266_), .B2(new_n274_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(new_n248_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n288_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT89), .A3(new_n274_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n286_), .A2(new_n287_), .B1(new_n248_), .B2(new_n290_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n274_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n299_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n293_), .B(new_n298_), .C1(new_n307_), .C2(new_n278_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G155gat), .B(G162gat), .Z(new_n309_));
  OR2_X1    g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n310_), .A2(KEYINPUT3), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(KEYINPUT3), .B2(new_n310_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT83), .Z(new_n316_));
  OAI21_X1  g115(.A(new_n309_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n309_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n310_), .A3(new_n312_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323_));
  XOR2_X1   g122(.A(G127gat), .B(G134gat), .Z(new_n324_));
  XOR2_X1   g123(.A(G113gat), .B(G120gat), .Z(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT90), .ZN(new_n329_));
  INV_X1    g128(.A(new_n322_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n322_), .A2(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n327_), .B(new_n329_), .C1(new_n334_), .C2(new_n323_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n332_), .A2(new_n333_), .A3(new_n328_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n291_), .B2(new_n284_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n278_), .B1(new_n275_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n307_), .B2(new_n278_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n308_), .B(new_n346_), .C1(new_n350_), .C2(new_n298_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n293_), .B1(new_n307_), .B2(new_n278_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n297_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n297_), .B(new_n293_), .C1(new_n307_), .C2(new_n278_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n327_), .B(new_n328_), .C1(new_n334_), .C2(new_n323_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n332_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n358_), .A2(KEYINPUT91), .A3(new_n339_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT91), .B1(new_n358_), .B2(new_n339_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT92), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n342_), .B(KEYINPUT33), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n351_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n305_), .B1(new_n322_), .B2(KEYINPUT29), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n330_), .B2(new_n368_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n322_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n366_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G228gat), .ZN(new_n374_));
  INV_X1    g173(.A(G233gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT84), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(KEYINPUT84), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n374_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G78gat), .ZN(new_n379_));
  INV_X1    g178(.A(G106gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n373_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(G43gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n249_), .A2(new_n265_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n249_), .B2(new_n265_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n326_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n391_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(new_n331_), .A3(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(G15gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT31), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n365_), .A2(new_n384_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n356_), .A2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n373_), .B(new_n383_), .Z(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n384_), .A3(new_n400_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n346_), .A2(KEYINPUT93), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n355_), .B(KEYINPUT27), .C1(new_n350_), .C2(new_n297_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n407_), .A2(new_n412_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n235_), .B1(new_n405_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G232gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT34), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n380_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G99gat), .A2(G106gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT6), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G99gat), .A3(G106gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT66), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G85gat), .A2(G92gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G85gat), .B(G92gat), .Z(new_n440_));
  AND2_X1   g239(.A1(new_n428_), .A2(new_n430_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  INV_X1    g241(.A(G99gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n380_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n440_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT8), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n431_), .A2(new_n445_), .A3(new_n444_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n440_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n439_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n423_), .B1(new_n452_), .B2(new_n211_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n449_), .A2(new_n450_), .A3(new_n440_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n449_), .B2(new_n440_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n448_), .A2(KEYINPUT68), .A3(new_n451_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n439_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n220_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n453_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n420_), .A2(new_n422_), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT72), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G190gat), .B(G218gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G134gat), .B(G162gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n468_), .A2(KEYINPUT36), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n453_), .B(new_n463_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n472_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n465_), .A2(new_n470_), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n468_), .B(KEYINPUT36), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT37), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n475_), .A2(KEYINPUT74), .A3(new_n476_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n471_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n487_));
  INV_X1    g286(.A(G71gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT67), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G71gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G78gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT67), .B(G71gat), .ZN(new_n494_));
  INV_X1    g293(.A(G78gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G64gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G57gat), .ZN(new_n499_));
  INV_X1    g298(.A(G57gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G64gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT11), .B1(new_n499_), .B2(new_n501_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n493_), .B(new_n496_), .C1(new_n502_), .C2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n487_), .B1(new_n452_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT64), .Z(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n452_), .B2(new_n507_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n506_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT12), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n508_), .B(new_n511_), .C1(new_n459_), .C2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n452_), .A2(new_n507_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n438_), .A2(new_n434_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n432_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(new_n512_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n510_), .B1(new_n515_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G120gat), .B(G148gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT5), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G176gat), .B(G204gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n514_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT70), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n514_), .A2(new_n521_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n525_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n528_), .A2(KEYINPUT13), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT13), .B1(new_n528_), .B2(new_n530_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n208_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(new_n507_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G127gat), .B(G155gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT16), .ZN(new_n540_));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n538_), .A2(new_n544_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n486_), .A2(new_n534_), .A3(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n418_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n415_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n203_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT38), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n481_), .A2(new_n471_), .A3(new_n483_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n405_), .B2(new_n417_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n534_), .A2(new_n235_), .A3(new_n548_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(G1gat), .B1(new_n560_), .B2(new_n415_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n552_), .A2(new_n553_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n554_), .A2(new_n561_), .A3(new_n562_), .ZN(G1324gat));
  NAND2_X1  g362(.A1(new_n407_), .A2(new_n416_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G8gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT39), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n550_), .A2(new_n204_), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT40), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(G1325gat));
  AOI21_X1  g370(.A(new_n396_), .B1(new_n559_), .B2(new_n403_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT41), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n550_), .A2(new_n396_), .A3(new_n403_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(G1326gat));
  NOR2_X1   g374(.A1(new_n384_), .A2(G22gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT95), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n550_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G22gat), .B1(new_n560_), .B2(new_n384_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT94), .B(KEYINPUT42), .Z(new_n580_));
  AND2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT96), .ZN(G1327gat));
  NAND2_X1  g383(.A1(new_n556_), .A2(new_n548_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n534_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n418_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G29gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n551_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n548_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n534_), .A2(new_n235_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT43), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n405_), .A2(new_n417_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(new_n486_), .ZN(new_n596_));
  AOI211_X1 g395(.A(KEYINPUT43), .B(new_n485_), .C1(new_n405_), .C2(new_n417_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT44), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT44), .B(new_n593_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n600_), .A2(new_n551_), .A3(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n591_), .B1(new_n602_), .B2(new_n590_), .ZN(G1328gat));
  AOI21_X1  g402(.A(G36gat), .B1(new_n407_), .B2(new_n416_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n589_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT45), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT45), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n589_), .A2(new_n607_), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n600_), .A2(new_n564_), .A3(new_n601_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT98), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n600_), .A2(KEYINPUT98), .A3(new_n564_), .A4(new_n601_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G36gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT46), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  OAI221_X1 g416(.A(new_n609_), .B1(new_n615_), .B2(KEYINPUT46), .C1(new_n611_), .C2(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1329gat));
  INV_X1    g418(.A(G43gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n589_), .A2(new_n620_), .A3(new_n403_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n600_), .A2(new_n403_), .A3(new_n601_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n622_), .B2(new_n620_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g423(.A(G50gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n589_), .A2(new_n625_), .A3(new_n408_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n600_), .A2(new_n408_), .A3(new_n601_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n628_), .A3(G50gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(G50gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(G1331gat));
  NAND2_X1  g430(.A1(new_n595_), .A2(new_n235_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n533_), .B1(new_n632_), .B2(KEYINPUT101), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(KEYINPUT101), .B2(new_n632_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(new_n548_), .A3(new_n486_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n500_), .A3(new_n551_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n557_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n534_), .A2(new_n235_), .A3(new_n592_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G57gat), .B1(new_n640_), .B2(new_n415_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(G1332gat));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n498_), .A3(new_n564_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n498_), .B1(new_n639_), .B2(new_n564_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT102), .B(KEYINPUT48), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n643_), .A2(new_n646_), .ZN(G1333gat));
  AOI21_X1  g446(.A(new_n488_), .B1(new_n639_), .B2(new_n403_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT49), .Z(new_n649_));
  NAND3_X1  g448(.A1(new_n635_), .A2(new_n488_), .A3(new_n403_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1334gat));
  AOI21_X1  g450(.A(new_n495_), .B1(new_n639_), .B2(new_n408_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT50), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n635_), .A2(new_n495_), .A3(new_n408_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1335gat));
  NOR2_X1   g454(.A1(new_n634_), .A2(new_n585_), .ZN(new_n656_));
  INV_X1    g455(.A(G85gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n551_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n534_), .A2(new_n235_), .A3(new_n548_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT103), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n661_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(KEYINPUT104), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n415_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n658_), .B1(new_n667_), .B2(new_n657_), .ZN(G1336gat));
  INV_X1    g467(.A(G92gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n656_), .A2(new_n669_), .A3(new_n564_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n665_), .A2(new_n666_), .B1(new_n407_), .B2(new_n416_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n669_), .ZN(G1337gat));
  OR2_X1    g471(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n665_), .A2(new_n666_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n403_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G99gat), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n403_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n656_), .A2(new_n677_), .B1(KEYINPUT105), .B2(KEYINPUT51), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n673_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n404_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n678_), .B(new_n673_), .C1(new_n680_), .C2(new_n443_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n679_), .A2(new_n682_), .ZN(G1338gat));
  XNOR2_X1  g482(.A(KEYINPUT107), .B(KEYINPUT53), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n408_), .B(new_n661_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G106gat), .B1(new_n685_), .B2(new_n686_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT52), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n685_), .A2(new_n686_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT52), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n687_), .A4(G106gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  NOR4_X1   g493(.A1(new_n634_), .A2(G106gat), .A3(new_n384_), .A4(new_n585_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n684_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n684_), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n695_), .B(new_n698_), .C1(new_n690_), .C2(new_n693_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1339gat));
  AND2_X1   g499(.A1(new_n234_), .A2(new_n528_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n452_), .A2(new_n507_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n508_), .B(new_n703_), .C1(new_n459_), .C2(new_n513_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n514_), .A2(KEYINPUT55), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n455_), .A2(new_n456_), .A3(new_n454_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT68), .B1(new_n448_), .B2(new_n451_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n518_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n513_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT55), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n508_), .A4(new_n511_), .ZN(new_n712_));
  AOI221_X4 g511(.A(new_n702_), .B1(new_n510_), .B2(new_n704_), .C1(new_n705_), .C2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n705_), .A2(new_n712_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n704_), .A2(new_n510_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT109), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n525_), .B1(new_n713_), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT110), .B(KEYINPUT56), .Z(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n717_), .A2(KEYINPUT111), .A3(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT56), .B(new_n525_), .C1(new_n713_), .C2(new_n716_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT111), .B1(new_n717_), .B2(new_n719_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n701_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n216_), .A2(new_n222_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n221_), .A2(new_n213_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(new_n231_), .C1(new_n726_), .C2(new_n222_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(new_n233_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n528_), .A2(new_n530_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n731_), .A2(KEYINPUT57), .A3(new_n555_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT57), .ZN(new_n733_));
  INV_X1    g532(.A(new_n730_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735_));
  INV_X1    g534(.A(new_n487_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n519_), .B2(new_n512_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n711_), .B1(new_n738_), .B2(new_n511_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n514_), .A2(KEYINPUT55), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n715_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n702_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n714_), .A2(KEYINPUT109), .A3(new_n715_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n526_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n735_), .B1(new_n744_), .B2(new_n718_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n721_), .A3(new_n720_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n734_), .B1(new_n746_), .B2(new_n701_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n733_), .B1(new_n747_), .B2(new_n556_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n728_), .A2(new_n528_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n717_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n752_), .B2(new_n721_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(KEYINPUT58), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n754_), .B2(new_n486_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n749_), .B(new_n486_), .C1(new_n753_), .C2(KEYINPUT58), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n752_), .A2(new_n721_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n728_), .A2(new_n528_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(KEYINPUT58), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT113), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n753_), .A2(new_n761_), .A3(KEYINPUT58), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n756_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n732_), .B(new_n748_), .C1(new_n755_), .C2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n548_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n486_), .A2(new_n548_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n235_), .A4(new_n533_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n549_), .A2(KEYINPUT108), .A3(new_n767_), .A4(new_n235_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n766_), .A2(new_n235_), .A3(new_n533_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT54), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n771_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n765_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n551_), .A2(new_n407_), .A3(new_n416_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n411_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(G113gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n234_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n764_), .A2(new_n782_), .A3(new_n548_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n764_), .B2(new_n548_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n774_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT59), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n770_), .A2(new_n773_), .A3(new_n771_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n548_), .B2(new_n764_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n777_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT59), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n234_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n781_), .B1(new_n795_), .B2(new_n780_), .ZN(G1340gat));
  XOR2_X1   g595(.A(KEYINPUT116), .B(G120gat), .Z(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n533_), .B2(KEYINPUT60), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n779_), .B(new_n798_), .C1(KEYINPUT60), .C2(new_n797_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n797_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n765_), .A2(KEYINPUT115), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n764_), .A2(new_n782_), .A3(new_n548_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n790_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n787_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n793_), .B(new_n534_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n800_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n533_), .B1(new_n778_), .B2(KEYINPUT59), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT117), .B1(new_n789_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n799_), .B1(new_n807_), .B2(new_n809_), .ZN(G1341gat));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n779_), .A2(new_n811_), .A3(new_n592_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n789_), .A2(new_n592_), .A3(new_n793_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n814_), .B2(new_n811_), .ZN(G1342gat));
  NAND4_X1  g614(.A1(new_n789_), .A2(G134gat), .A3(new_n486_), .A4(new_n793_), .ZN(new_n816_));
  INV_X1    g615(.A(G134gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n778_), .B2(new_n555_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n819_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n816_), .A2(new_n820_), .A3(new_n821_), .ZN(G1343gat));
  NOR2_X1   g621(.A1(new_n776_), .A2(new_n409_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n775_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n234_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n534_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g628(.A1(new_n824_), .A2(new_n548_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT61), .B(G155gat), .Z(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1346gat));
  INV_X1    g631(.A(G162gat), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n824_), .A2(new_n833_), .A3(new_n485_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n824_), .B2(new_n555_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n836_), .B2(new_n837_), .ZN(G1347gat));
  INV_X1    g637(.A(KEYINPUT22), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n551_), .B1(new_n407_), .B2(new_n416_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n403_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT120), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n843_), .A3(new_n403_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n408_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n785_), .A2(new_n839_), .A3(new_n234_), .A4(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n848_), .A2(KEYINPUT62), .A3(new_n250_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT62), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n785_), .A2(new_n851_), .A3(new_n234_), .A4(new_n847_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n852_), .A2(G169gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n850_), .B2(new_n853_), .ZN(G1348gat));
  AND2_X1   g653(.A1(new_n785_), .A2(new_n847_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G176gat), .B1(new_n855_), .B2(new_n534_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n791_), .A2(new_n408_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n846_), .A2(new_n251_), .A3(new_n533_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1349gat));
  NOR2_X1   g658(.A1(new_n548_), .A2(new_n279_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n785_), .A2(new_n847_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n862_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n846_), .A2(new_n548_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G183gat), .B1(new_n857_), .B2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n863_), .A2(new_n864_), .A3(new_n866_), .ZN(G1350gat));
  NAND4_X1  g666(.A1(new_n855_), .A2(new_n259_), .A3(new_n263_), .A4(new_n556_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n785_), .A2(new_n486_), .A3(new_n847_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n869_), .A2(new_n870_), .A3(G190gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(G190gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(G1351gat));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n840_), .A2(new_n408_), .A3(new_n404_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n791_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n775_), .A2(KEYINPUT123), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n234_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g680(.A(new_n533_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n882_));
  INV_X1    g681(.A(G204gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(KEYINPUT124), .B2(new_n883_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT124), .B(G204gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n882_), .B2(new_n885_), .ZN(G1353gat));
  AOI21_X1  g685(.A(new_n548_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT125), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1354gat));
  NAND2_X1  g690(.A1(new_n879_), .A2(new_n556_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n555_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G218gat), .B1(new_n895_), .B2(KEYINPUT126), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n486_), .A2(G218gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT127), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n894_), .A2(new_n896_), .B1(new_n879_), .B2(new_n898_), .ZN(G1355gat));
endmodule


