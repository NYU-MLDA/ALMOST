//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_;
  INV_X1    g000(.A(G197gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G197gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT21), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT91), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT92), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT92), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT90), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n203_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n202_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n205_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT21), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n208_), .A2(new_n212_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n209_), .B(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n206_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n224_), .B(KEYINPUT87), .Z(new_n225_));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(KEYINPUT1), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n229_), .B(KEYINPUT3), .Z(new_n233_));
  XOR2_X1   g032(.A(new_n231_), .B(KEYINPUT2), .Z(new_n234_));
  OAI211_X1 g033(.A(new_n225_), .B(new_n226_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n223_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G22gat), .B(G50gat), .Z(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  AND2_X1   g039(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(G233gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(G78gat), .Z(new_n244_));
  INV_X1    g043(.A(G106gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n232_), .A2(new_n235_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n250_), .A2(KEYINPUT29), .A3(new_n247_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n246_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n240_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n240_), .B1(new_n253_), .B2(new_n252_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT27), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G226gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT19), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT76), .ZN(new_n262_));
  INV_X1    g061(.A(G183gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT25), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n263_), .A2(KEYINPUT25), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n261_), .B(new_n264_), .C1(new_n265_), .C2(new_n262_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT77), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT24), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT23), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G183gat), .A3(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n269_), .A2(KEYINPUT24), .A3(new_n279_), .A4(new_n270_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n266_), .A2(new_n273_), .A3(new_n278_), .A4(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT79), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n277_), .A2(KEYINPUT79), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n290_), .B2(G169gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n288_), .B(new_n291_), .C1(new_n292_), .C2(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n279_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n281_), .B1(new_n287_), .B2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n295_), .C2(new_n223_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT25), .B(G183gat), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n261_), .A2(new_n297_), .B1(new_n272_), .B2(new_n267_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n283_), .A2(new_n298_), .A3(new_n286_), .A4(new_n280_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n292_), .A2(new_n288_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n300_), .B(new_n279_), .C1(new_n282_), .C2(new_n284_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n210_), .A2(new_n211_), .B1(new_n216_), .B2(KEYINPUT21), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n303_), .A2(new_n208_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n296_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n279_), .A3(new_n293_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n308_), .A3(new_n281_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT93), .B1(new_n309_), .B2(KEYINPUT20), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n260_), .B1(new_n306_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT20), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n260_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n295_), .A2(new_n223_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT95), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT94), .B(KEYINPUT18), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  AND3_X1   g121(.A1(new_n311_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n258_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n311_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT99), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n315_), .B1(new_n313_), .B2(new_n327_), .ZN(new_n328_));
  AOI211_X1 g127(.A(KEYINPUT99), .B(new_n312_), .C1(new_n302_), .C2(new_n304_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n260_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT20), .B1(new_n295_), .B2(new_n223_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n333_), .A2(new_n314_), .A3(new_n305_), .A4(new_n296_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT27), .B(new_n326_), .C1(new_n335_), .C2(new_n322_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n325_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G120gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G113gat), .ZN(new_n339_));
  INV_X1    g138(.A(G113gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G120gat), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT82), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT82), .B1(new_n339_), .B2(new_n341_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G127gat), .B(G134gat), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G127gat), .B(G134gat), .Z(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n340_), .A2(G120gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n338_), .A2(G113gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n339_), .A2(new_n341_), .A3(KEYINPUT82), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n353_), .A2(KEYINPUT83), .A3(KEYINPUT84), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n344_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n355_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n346_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT84), .B1(new_n353_), .B2(KEYINPUT83), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n357_), .A3(new_n355_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n345_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n364_), .B(G15gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(G71gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT80), .B(G43gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G99gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n366_), .B(new_n368_), .Z(new_n369_));
  NAND3_X1  g168(.A1(new_n308_), .A2(KEYINPUT30), .A3(new_n281_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT30), .B1(new_n308_), .B2(new_n281_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT81), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n295_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n370_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n369_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n369_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT31), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n369_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n371_), .A2(new_n372_), .A3(KEYINPUT81), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n376_), .B1(new_n375_), .B2(new_n370_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT31), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n379_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n381_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n381_), .B2(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n363_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n381_), .A2(new_n387_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT85), .ZN(new_n393_));
  INV_X1    g192(.A(new_n363_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n381_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AND4_X1   g195(.A1(new_n257_), .A2(new_n337_), .A3(new_n391_), .A4(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n359_), .A2(new_n362_), .A3(new_n250_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n232_), .B(new_n235_), .C1(new_n345_), .C2(new_n353_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(KEYINPUT4), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n398_), .A2(KEYINPUT96), .A3(KEYINPUT4), .A4(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n359_), .A2(new_n405_), .A3(new_n362_), .A4(new_n250_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n404_), .A2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n398_), .A2(new_n399_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n407_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G85gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  NAND3_X1  g216(.A1(new_n411_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n417_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n409_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n413_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n397_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n256_), .A2(new_n336_), .A3(new_n325_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(new_n423_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n311_), .A2(new_n316_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(new_n330_), .B2(new_n334_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n417_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n420_), .A2(new_n421_), .A3(new_n419_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT100), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n406_), .A2(new_n407_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n404_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT98), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n398_), .A2(new_n399_), .A3(new_n408_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n419_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT97), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT98), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n404_), .A2(new_n444_), .A3(new_n437_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n418_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n323_), .A2(new_n324_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n411_), .A2(KEYINPUT33), .A3(new_n413_), .A4(new_n417_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n446_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n423_), .A2(KEYINPUT100), .A3(new_n431_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n436_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n427_), .B1(new_n453_), .B2(new_n257_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n391_), .A2(new_n396_), .A3(KEYINPUT86), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT86), .B1(new_n391_), .B2(new_n396_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n425_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT72), .B(G15gat), .ZN(new_n459_));
  INV_X1    g258(.A(G22gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G1gat), .B(G8gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n467_), .B(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n467_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n470_), .B(KEYINPUT15), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n467_), .A2(new_n470_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n472_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G113gat), .B(G141gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT74), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n474_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT75), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n458_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n494_));
  XOR2_X1   g293(.A(G71gat), .B(G78gat), .Z(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n494_), .A2(new_n495_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G231gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT73), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n475_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n503_));
  XOR2_X1   g302(.A(G127gat), .B(G155gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT16), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G183gat), .B(G211gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  OR3_X1    g306(.A1(new_n502_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(KEYINPUT17), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT6), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT64), .B(G85gat), .Z(new_n515_));
  INV_X1    g314(.A(KEYINPUT9), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(G92gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(G85gat), .B(G92gat), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT10), .B(G99gat), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n245_), .ZN(new_n521_));
  AND4_X1   g320(.A1(new_n514_), .A2(new_n517_), .A3(new_n519_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G85gat), .B(G92gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT7), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n526_), .B2(new_n514_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(KEYINPUT65), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n523_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT65), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n526_), .A2(new_n514_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(new_n524_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(KEYINPUT65), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT8), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n535_), .A2(new_n476_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n534_), .A3(new_n470_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT34), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(KEYINPUT67), .A3(new_n542_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n540_), .A2(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n547_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT68), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT69), .B(KEYINPUT36), .Z(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n512_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n553_), .B(KEYINPUT70), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT36), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n558_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n548_), .A2(new_n549_), .ZN(new_n564_));
  OAI221_X1 g363(.A(new_n556_), .B1(new_n557_), .B2(new_n512_), .C1(new_n564_), .C2(new_n561_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n511_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n498_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n535_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n529_), .A2(new_n534_), .A3(new_n498_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT12), .ZN(new_n573_));
  AOI211_X1 g372(.A(new_n573_), .B(new_n498_), .C1(new_n529_), .C2(new_n534_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n535_), .A2(KEYINPUT12), .A3(new_n569_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(KEYINPUT66), .A3(new_n571_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT12), .B1(new_n535_), .B2(new_n569_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n576_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n572_), .B1(new_n580_), .B2(new_n568_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G120gat), .B(G148gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n586_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n567_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n491_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n423_), .B(KEYINPUT101), .Z(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(G1gat), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n595_), .A2(new_n597_), .B1(KEYINPUT103), .B2(KEYINPUT38), .ZN(new_n598_));
  NOR2_X1   g397(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  NOR2_X1   g399(.A1(new_n559_), .A2(new_n562_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n458_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n488_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n593_), .A2(new_n511_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n424_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT102), .Z(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(KEYINPUT40), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n611_));
  INV_X1    g410(.A(new_n337_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n603_), .A2(new_n612_), .A3(new_n605_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(G8gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(G8gat), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(KEYINPUT105), .A3(new_n615_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n618_), .A2(new_n620_), .A3(KEYINPUT39), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n595_), .A2(new_n463_), .A3(new_n612_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n618_), .B2(KEYINPUT39), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n610_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n618_), .A2(KEYINPUT39), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n620_), .A3(KEYINPUT39), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(KEYINPUT40), .A3(new_n626_), .A4(new_n622_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(new_n457_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G15gat), .B1(new_n606_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  INV_X1    g430(.A(new_n595_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(G15gat), .A3(new_n629_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1326gat));
  OAI21_X1  g433(.A(G22gat), .B1(new_n606_), .B2(new_n257_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n595_), .A2(new_n460_), .A3(new_n256_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1327gat));
  INV_X1    g437(.A(new_n511_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n593_), .A2(new_n639_), .A3(new_n604_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n563_), .A2(new_n565_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n458_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n641_), .B1(new_n458_), .B2(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT44), .B(new_n640_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(G29gat), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n596_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n511_), .A2(new_n601_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n593_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n491_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n491_), .A2(KEYINPUT106), .A3(new_n653_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n423_), .A3(new_n657_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n649_), .A2(new_n651_), .B1(new_n650_), .B2(new_n658_), .ZN(G1328gat));
  NOR2_X1   g458(.A1(new_n337_), .A2(G36gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n657_), .A3(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n647_), .A2(new_n612_), .A3(new_n648_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT107), .B1(new_n664_), .B2(G36gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI221_X1 g468(.A(new_n663_), .B1(KEYINPUT109), .B2(KEYINPUT46), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  NAND2_X1  g470(.A1(new_n391_), .A2(new_n396_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n649_), .A2(G43gat), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n457_), .A3(new_n657_), .ZN(new_n675_));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g478(.A(G50gat), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n257_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n656_), .A2(new_n256_), .A3(new_n657_), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n649_), .A2(new_n681_), .B1(new_n680_), .B2(new_n682_), .ZN(G1331gat));
  INV_X1    g482(.A(new_n593_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n684_), .A2(new_n511_), .A3(new_n490_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n603_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G57gat), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n424_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n458_), .A2(new_n604_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n684_), .A2(new_n567_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n596_), .B1(new_n691_), .B2(KEYINPUT110), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(KEYINPUT110), .B2(new_n691_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n688_), .B1(new_n693_), .B2(new_n687_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n686_), .B2(new_n337_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT48), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT48), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n337_), .A2(G64gat), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT111), .ZN(new_n699_));
  OAI22_X1  g498(.A1(new_n696_), .A2(new_n697_), .B1(new_n691_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n686_), .B2(new_n629_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n629_), .A2(G71gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n691_), .B2(new_n704_), .ZN(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n686_), .B2(new_n257_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n257_), .A2(G78gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n707_), .B1(new_n691_), .B2(new_n708_), .ZN(G1335gat));
  AND4_X1   g508(.A1(new_n601_), .A2(new_n689_), .A3(new_n511_), .A4(new_n593_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n596_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G85gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n643_), .A2(new_n644_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n684_), .A2(new_n639_), .A3(new_n488_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT113), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n423_), .A2(new_n515_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT114), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n712_), .B1(new_n716_), .B2(new_n718_), .ZN(G1336gat));
  AOI21_X1  g518(.A(G92gat), .B1(new_n710_), .B2(new_n612_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT115), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n612_), .A2(G92gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n716_), .B2(new_n722_), .ZN(G1337gat));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n457_), .A3(new_n714_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n673_), .A2(new_n520_), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n724_), .A2(G99gat), .B1(new_n710_), .B2(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n245_), .A3(new_n256_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n256_), .A3(new_n714_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n733_), .B(new_n735_), .ZN(G1339gat));
  INV_X1    g535(.A(KEYINPUT120), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT57), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n588_), .A2(new_n488_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n570_), .A2(new_n573_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(KEYINPUT66), .A3(new_n571_), .A4(new_n577_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n568_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n576_), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT55), .B(new_n742_), .C1(new_n741_), .C2(new_n576_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n580_), .B2(new_n568_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n585_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n739_), .B1(new_n748_), .B2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n747_), .A2(new_n749_), .A3(new_n750_), .A4(new_n585_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n471_), .A2(new_n472_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n477_), .A2(new_n478_), .A3(new_n473_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n485_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n487_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n752_), .A2(new_n753_), .B1(new_n589_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n738_), .B1(new_n759_), .B2(new_n601_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n748_), .A2(new_n751_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n739_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n753_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n589_), .A2(new_n758_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT57), .A3(new_n602_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n743_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n577_), .A2(KEYINPUT66), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n571_), .A2(KEYINPUT66), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n574_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n770_), .B2(new_n740_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT55), .B1(new_n771_), .B2(new_n742_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n580_), .A2(new_n745_), .A3(new_n568_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n767_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n586_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n747_), .A2(new_n750_), .A3(new_n585_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n588_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n757_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT58), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .A4(KEYINPUT58), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n642_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n760_), .A2(new_n766_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n511_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n566_), .A2(new_n592_), .A3(new_n591_), .A4(new_n489_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT54), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n684_), .A2(new_n788_), .A3(new_n489_), .A4(new_n566_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n785_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n711_), .A2(new_n397_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n489_), .A2(new_n340_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n790_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n783_), .A2(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n781_), .A2(new_n800_), .A3(new_n642_), .A4(new_n782_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n799_), .A2(new_n801_), .A3(new_n760_), .A4(new_n766_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n798_), .B1(new_n802_), .B2(new_n511_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT59), .B1(new_n803_), .B2(new_n792_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n803_), .C2(new_n792_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n795_), .B(new_n797_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n803_), .A2(new_n792_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n488_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n737_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n806_), .A2(new_n807_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(KEYINPUT120), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(G1340gat));
  XNOR2_X1  g615(.A(KEYINPUT121), .B(G120gat), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n593_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n809_), .B1(KEYINPUT60), .B2(new_n818_), .ZN(new_n819_));
  AND4_X1   g618(.A1(new_n593_), .A2(new_n812_), .A3(new_n794_), .A4(new_n819_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n820_), .A2(new_n817_), .B1(KEYINPUT60), .B2(new_n819_), .ZN(G1341gat));
  INV_X1    g620(.A(G127gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n809_), .A2(new_n822_), .A3(new_n639_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n511_), .B(new_n795_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n822_), .ZN(G1342gat));
  INV_X1    g624(.A(G134gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n809_), .A2(new_n826_), .A3(new_n601_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n642_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n795_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n829_), .B2(new_n826_), .ZN(G1343gat));
  INV_X1    g629(.A(new_n803_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n457_), .A2(new_n426_), .A3(new_n596_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n488_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g635(.A1(new_n833_), .A2(new_n684_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT122), .B(G148gat), .Z(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1345gat));
  NOR2_X1   g638(.A1(new_n833_), .A2(new_n511_), .ZN(new_n840_));
  XOR2_X1   g639(.A(KEYINPUT61), .B(G155gat), .Z(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1346gat));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n834_), .B2(new_n642_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n833_), .A2(G162gat), .A3(new_n602_), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n844_), .B2(new_n846_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1347gat));
  NAND2_X1  g648(.A1(new_n791_), .A2(new_n257_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n629_), .A2(new_n337_), .A3(new_n711_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n292_), .A3(new_n488_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n850_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n488_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT124), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n858_), .A2(new_n859_), .A3(G169gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n858_), .B2(G169gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n854_), .B1(new_n860_), .B2(new_n861_), .ZN(G1348gat));
  AOI21_X1  g661(.A(G176gat), .B1(new_n853_), .B2(new_n593_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n803_), .A2(new_n256_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n852_), .A2(new_n288_), .A3(new_n684_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1349gat));
  NAND2_X1  g665(.A1(new_n851_), .A2(new_n639_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n850_), .A2(new_n297_), .A3(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT125), .ZN(new_n869_));
  INV_X1    g668(.A(new_n867_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G183gat), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1350gat));
  NAND3_X1  g671(.A1(new_n853_), .A2(new_n261_), .A3(new_n601_), .ZN(new_n873_));
  INV_X1    g672(.A(G190gat), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n850_), .A2(new_n828_), .A3(new_n852_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1351gat));
  NOR4_X1   g675(.A1(new_n457_), .A2(new_n423_), .A3(new_n257_), .A4(new_n337_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n831_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n604_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n202_), .ZN(G1352gat));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n684_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n204_), .ZN(G1353gat));
  INV_X1    g681(.A(new_n878_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n884_));
  INV_X1    g683(.A(G211gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n639_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT126), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n885_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1354gat));
  AND3_X1   g689(.A1(new_n883_), .A2(G218gat), .A3(new_n642_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n878_), .A2(new_n602_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT127), .ZN(new_n893_));
  AOI21_X1  g692(.A(G218gat), .B1(new_n892_), .B2(KEYINPUT127), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(G1355gat));
endmodule


