//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT84), .B(KEYINPUT2), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n202_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(KEYINPUT84), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(KEYINPUT84), .ZN(new_n209_));
  OAI211_X1 g008(.A(KEYINPUT85), .B(new_n204_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT3), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n212_), .A2(new_n214_), .B1(new_n205_), .B2(KEYINPUT2), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n206_), .A2(new_n210_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT83), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n219_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n205_), .A2(new_n211_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G127gat), .B(G134gat), .Z(new_n231_));
  XOR2_X1   g030(.A(G113gat), .B(G120gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n216_), .A2(new_n220_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G1gat), .B(G29gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n238_), .B(KEYINPUT93), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n221_), .A2(new_n233_), .A3(new_n229_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n233_), .B1(new_n221_), .B2(new_n229_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n247_), .B1(new_n250_), .B2(KEYINPUT4), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n230_), .A2(new_n252_), .A3(new_n234_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT94), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n249_), .A2(KEYINPUT94), .A3(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n245_), .B1(new_n251_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT96), .B1(new_n258_), .B2(KEYINPUT33), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n235_), .A2(KEYINPUT4), .A3(new_n237_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT94), .B1(new_n249_), .B2(new_n252_), .ZN(new_n261_));
  NOR4_X1   g060(.A1(new_n236_), .A2(new_n254_), .A3(KEYINPUT4), .A4(new_n233_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n260_), .B(new_n246_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n244_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n250_), .B2(new_n238_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT96), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n260_), .B(new_n238_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT97), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT97), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n257_), .A2(new_n272_), .A3(new_n260_), .A4(new_n238_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n235_), .A2(new_n237_), .A3(new_n246_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n264_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(new_n269_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n258_), .A2(KEYINPUT33), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n283_), .B(new_n284_), .C1(G183gat), .C2(G190gat), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT79), .B1(new_n286_), .B2(KEYINPUT22), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT22), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(G169gat), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT78), .B1(new_n289_), .B2(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n286_), .A3(KEYINPUT22), .ZN(new_n294_));
  INV_X1    g093(.A(G176gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n280_), .B(new_n285_), .C1(new_n291_), .C2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT26), .B(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G183gat), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(new_n299_), .B2(G183gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n298_), .A2(new_n300_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n283_), .A2(new_n284_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(G169gat), .B2(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n286_), .A2(new_n295_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n305_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n297_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G197gat), .A2(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT21), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(KEYINPUT21), .A3(new_n316_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n289_), .A2(G169gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n286_), .A2(KEYINPUT22), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n295_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n285_), .A2(new_n280_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT25), .B(G183gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n298_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n312_), .A2(new_n332_), .A3(new_n307_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT90), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n306_), .B1(new_n298_), .B2(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n312_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n330_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n325_), .B(KEYINPUT20), .C1(new_n338_), .C2(new_n324_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT91), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n338_), .B2(new_n324_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT20), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n297_), .A2(new_n313_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n322_), .A2(new_n323_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n343_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n336_), .B1(new_n335_), .B2(new_n312_), .ZN(new_n350_));
  AND4_X1   g149(.A1(new_n336_), .A2(new_n312_), .A3(new_n332_), .A4(new_n307_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n324_), .B(new_n329_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n341_), .ZN(new_n353_));
  AND4_X1   g152(.A1(new_n343_), .A2(new_n352_), .A3(new_n348_), .A4(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n342_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n342_), .B(new_n360_), .C1(new_n349_), .C2(new_n354_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n279_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n244_), .B1(new_n263_), .B2(new_n239_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n266_), .A2(KEYINPUT98), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT98), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n263_), .A2(new_n265_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n365_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n333_), .A2(new_n322_), .A3(new_n329_), .A4(new_n323_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT20), .B(new_n370_), .C1(new_n314_), .C2(new_n324_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n341_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n355_), .B2(new_n374_), .ZN(new_n376_));
  OAI22_X1  g175(.A1(new_n278_), .A2(new_n364_), .B1(new_n369_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT86), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n221_), .B2(new_n229_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n382_), .B2(new_n324_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n347_), .B(new_n379_), .C1(new_n236_), .C2(new_n381_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G78gat), .B(G106gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G22gat), .B(G50gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT28), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n236_), .A2(new_n389_), .A3(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n236_), .B2(new_n381_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(new_n390_), .A3(new_n387_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n383_), .A2(new_n384_), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n385_), .B(KEYINPUT87), .Z(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n399_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n397_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT88), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n383_), .A2(new_n384_), .A3(new_n402_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n403_), .A2(KEYINPUT88), .B1(new_n393_), .B2(new_n395_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n401_), .A2(new_n404_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT27), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n360_), .B(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n373_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n363_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT100), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT100), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n414_), .A2(new_n363_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n362_), .A2(new_n363_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n416_), .A2(new_n418_), .B1(new_n419_), .B2(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n263_), .A2(new_n239_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n264_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n263_), .A2(new_n265_), .A3(new_n367_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n367_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n410_), .A2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n377_), .A2(new_n410_), .B1(new_n420_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT80), .B(G15gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G227gat), .ZN(new_n430_));
  INV_X1    g229(.A(G233gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n297_), .A2(new_n313_), .A3(KEYINPUT30), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT30), .B1(new_n297_), .B2(new_n313_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n346_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n432_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n433_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441_));
  INV_X1    g240(.A(G43gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n436_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n429_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n428_), .A3(new_n445_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .A4(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n454_), .A2(new_n234_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n234_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT101), .B1(new_n427_), .B2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n362_), .A2(new_n363_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n414_), .A2(new_n417_), .A3(new_n363_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n417_), .B1(new_n414_), .B2(new_n363_), .ZN(new_n463_));
  OAI22_X1  g262(.A1(new_n461_), .A2(KEYINPUT27), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n396_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n400_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n404_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n408_), .A2(new_n409_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n464_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n459_), .A2(new_n369_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n454_), .A2(new_n456_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n233_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n454_), .A2(new_n234_), .A3(new_n456_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT101), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n266_), .A2(new_n268_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n275_), .B1(new_n270_), .B2(KEYINPUT97), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n477_), .A2(KEYINPUT96), .B1(new_n478_), .B2(new_n273_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n479_), .A2(new_n461_), .A3(new_n279_), .A4(new_n269_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n355_), .A2(new_n374_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n425_), .A2(new_n481_), .A3(new_n375_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n469_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n469_), .A2(new_n369_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n464_), .A2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n475_), .B(new_n476_), .C1(new_n483_), .C2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n460_), .A2(new_n471_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT74), .B(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G29gat), .B(G36gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n497_), .A2(new_n498_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n496_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n497_), .A2(new_n498_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT15), .A3(new_n499_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n495_), .A2(new_n502_), .A3(new_n503_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n499_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n503_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n493_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n511_), .B(KEYINPUT75), .Z(new_n512_));
  NAND3_X1  g311(.A1(new_n506_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT76), .ZN(new_n514_));
  INV_X1    g313(.A(new_n511_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n495_), .A2(new_n503_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(new_n507_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n507_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n495_), .B2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT76), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n506_), .A2(new_n510_), .A3(new_n521_), .A4(new_n512_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G169gat), .B(G197gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n514_), .A2(new_n520_), .A3(new_n522_), .A4(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n487_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G85gat), .B(G92gat), .Z(new_n532_));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI22_X1  g337(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n532_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT8), .B(new_n532_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n532_), .A2(KEYINPUT9), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT10), .B(G99gat), .Z(new_n546_));
  INV_X1    g345(.A(G106gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n533_), .B(KEYINPUT6), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT64), .B(G85gat), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT9), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(G92gat), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n545_), .A2(new_n548_), .A3(new_n549_), .A4(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n543_), .A2(new_n544_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(KEYINPUT12), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT66), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT66), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n554_), .A2(new_n564_), .A3(KEYINPUT12), .A4(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n554_), .A2(new_n561_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n554_), .A2(new_n561_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT12), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n568_), .ZN(new_n573_));
  OAI211_X1 g372(.A(G230gat), .B(G233gat), .C1(new_n573_), .C2(new_n569_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G120gat), .B(G148gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT67), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n575_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT13), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n561_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n516_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XOR2_X1   g389(.A(G183gat), .B(G211gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n587_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n554_), .A2(new_n518_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n554_), .A2(new_n505_), .A3(new_n502_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT70), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n598_), .A2(KEYINPUT71), .A3(new_n603_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n608_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .A4(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n601_), .A2(new_n602_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n604_), .A2(new_n607_), .A3(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT72), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n614_), .A2(new_n616_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n597_), .B1(new_n623_), .B2(KEYINPUT73), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n615_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n619_), .B(new_n620_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  OAI221_X1 g427(.A(new_n623_), .B1(KEYINPUT73), .B2(new_n597_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n596_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n531_), .A2(new_n584_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n488_), .A3(new_n425_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n487_), .A2(new_n627_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n530_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n583_), .A2(new_n636_), .A3(new_n596_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT102), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n369_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(new_n633_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n634_), .A2(new_n640_), .A3(new_n641_), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n631_), .A2(new_n489_), .A3(new_n464_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G8gat), .B1(new_n639_), .B2(new_n420_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1325gat));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n631_), .A2(new_n650_), .A3(new_n459_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G15gat), .B1(new_n639_), .B2(new_n475_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n639_), .B2(new_n410_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n410_), .A2(G22gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n631_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1327gat));
  NOR3_X1   g463(.A1(new_n583_), .A2(new_n595_), .A3(new_n627_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n531_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n425_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n583_), .A2(new_n636_), .A3(new_n595_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n628_), .A2(new_n629_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n487_), .A2(new_n669_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n487_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(KEYINPUT44), .B(new_n668_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n425_), .A2(G29gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n667_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  NOR2_X1   g479(.A1(new_n420_), .A2(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n531_), .A2(new_n665_), .A3(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n531_), .A2(new_n665_), .A3(new_n681_), .A4(new_n683_), .ZN(new_n686_));
  OR2_X1    g485(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n676_), .A2(new_n464_), .A3(new_n677_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G36gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT107), .Z(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n690_), .B(new_n693_), .ZN(G1329gat));
  NOR2_X1   g493(.A1(new_n475_), .A2(new_n442_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n676_), .A2(new_n677_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT108), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n676_), .A2(new_n698_), .A3(new_n677_), .A4(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n666_), .A2(new_n459_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n442_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n699_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT47), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n697_), .A2(new_n704_), .A3(new_n699_), .A4(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1330gat));
  AOI21_X1  g505(.A(G50gat), .B1(new_n666_), .B2(new_n469_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n469_), .A2(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n678_), .B2(new_n708_), .ZN(G1331gat));
  NAND2_X1  g508(.A1(new_n583_), .A2(new_n636_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(new_n596_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n635_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n369_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n487_), .A2(new_n636_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n715_), .A2(new_n583_), .A3(new_n630_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n425_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n720_), .A3(new_n464_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n712_), .A2(new_n464_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G64gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT110), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n725_), .A3(G64gat), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n724_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n721_), .B1(new_n728_), .B2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n712_), .B2(new_n459_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT49), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n716_), .A2(new_n731_), .A3(new_n459_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1334gat));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n712_), .B2(new_n469_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT50), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n716_), .A2(new_n736_), .A3(new_n469_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1335gat));
  INV_X1    g539(.A(new_n627_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n583_), .A2(new_n715_), .A3(new_n596_), .A4(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G85gat), .B1(new_n742_), .B2(new_n425_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n672_), .A2(new_n673_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n710_), .A2(new_n595_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n425_), .A2(new_n550_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  OAI21_X1  g548(.A(G92gat), .B1(new_n746_), .B2(new_n420_), .ZN(new_n750_));
  INV_X1    g549(.A(G92gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n742_), .A2(new_n751_), .A3(new_n464_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1337gat));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n754_));
  OAI21_X1  g553(.A(G99gat), .B1(new_n746_), .B2(new_n475_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n742_), .A2(new_n459_), .A3(new_n546_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n754_), .B(KEYINPUT51), .C1(new_n755_), .C2(new_n756_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n759_));
  AND4_X1   g558(.A1(new_n758_), .A2(new_n755_), .A3(new_n759_), .A4(new_n756_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n742_), .A2(new_n547_), .A3(new_n469_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n469_), .B(new_n745_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n512_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n506_), .A2(new_n510_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n770_), .B(new_n527_), .C1(new_n771_), .C2(new_n512_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n529_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n529_), .A2(new_n772_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT115), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n582_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n580_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n572_), .A2(new_n574_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n530_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT113), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n530_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n567_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n572_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n566_), .A2(KEYINPUT55), .A3(new_n567_), .A4(new_n571_), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n785_), .B(new_n778_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(KEYINPUT114), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n789_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n580_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n785_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(KEYINPUT56), .A3(new_n580_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n777_), .B1(new_n791_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n769_), .B1(new_n798_), .B2(new_n741_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n776_), .A2(new_n774_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n580_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n800_), .B(new_n779_), .C1(new_n801_), .C2(new_n790_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n803_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n671_), .A3(new_n805_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n801_), .A2(new_n790_), .A3(KEYINPUT114), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n783_), .B(new_n781_), .C1(new_n796_), .C2(new_n795_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n627_), .C1(new_n809_), .C2(new_n777_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n799_), .A2(new_n806_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n596_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n630_), .A2(new_n584_), .A3(new_n636_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n459_), .A2(new_n425_), .A3(new_n470_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT59), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n817_), .C1(new_n812_), .C2(new_n815_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n636_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n817_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n530_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n822_), .B2(new_n584_), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n584_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n824_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1341gat));
  XOR2_X1   g631(.A(KEYINPUT117), .B(G127gat), .Z(new_n833_));
  NOR2_X1   g632(.A1(new_n596_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT116), .B(G127gat), .C1(new_n824_), .C2(new_n595_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n816_), .A2(new_n595_), .A3(new_n818_), .ZN(new_n838_));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n836_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n835_), .B(KEYINPUT118), .C1(new_n836_), .C2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1342gat));
  XNOR2_X1  g644(.A(KEYINPUT119), .B(G134gat), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n822_), .A2(new_n670_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G134gat), .B1(new_n824_), .B2(new_n741_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1343gat));
  NAND4_X1  g648(.A1(new_n475_), .A2(new_n469_), .A3(new_n425_), .A4(new_n420_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n530_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n583_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n595_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  INV_X1    g657(.A(G162gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n851_), .A2(new_n859_), .A3(new_n741_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n851_), .A2(new_n671_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n859_), .ZN(G1347gat));
  AOI21_X1  g661(.A(new_n420_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n475_), .A2(new_n469_), .A3(new_n425_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865_), .B2(new_n636_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n865_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n869_), .A2(new_n530_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n867_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(new_n870_), .A3(new_n871_), .ZN(G1348gat));
  NOR2_X1   g671(.A1(new_n865_), .A2(new_n584_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n295_), .ZN(G1349gat));
  NOR2_X1   g673(.A1(new_n865_), .A2(new_n596_), .ZN(new_n875_));
  MUX2_X1   g674(.A(G183gat), .B(new_n331_), .S(new_n875_), .Z(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n865_), .B2(new_n670_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n741_), .A2(new_n298_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n865_), .B2(new_n878_), .ZN(G1351gat));
  NAND2_X1  g678(.A1(new_n475_), .A2(new_n426_), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT121), .Z(new_n881_));
  NAND2_X1  g680(.A1(new_n863_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n530_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(KEYINPUT122), .A2(G197gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(KEYINPUT122), .A2(G197gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT123), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1352gat));
  NOR2_X1   g689(.A1(new_n882_), .A2(new_n584_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G204gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n891_), .B(new_n893_), .ZN(G1353gat));
  NOR2_X1   g693(.A1(new_n882_), .A2(new_n596_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT63), .B(G211gat), .Z(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n895_), .B2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT126), .B(new_n902_), .C1(new_n882_), .C2(new_n596_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n898_), .A2(new_n900_), .B1(new_n904_), .B2(new_n905_), .ZN(G1354gat));
  XOR2_X1   g705(.A(KEYINPUT127), .B(G218gat), .Z(new_n907_));
  NOR3_X1   g706(.A1(new_n882_), .A2(new_n670_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n883_), .A2(new_n741_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1355gat));
endmodule


