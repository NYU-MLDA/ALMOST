//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XOR2_X1   g001(.A(G57gat), .B(G64gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n203_), .A2(new_n204_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT65), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  AND2_X1   g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G85gat), .B(G92gat), .Z(new_n222_));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT10), .B(G99gat), .Z(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n223_), .A2(new_n224_), .A3(G85gat), .A4(G92gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n221_), .A2(new_n227_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  OR3_X1    g032(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n222_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(new_n235_), .B2(new_n222_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n232_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n213_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT12), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(KEYINPUT66), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n232_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n213_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n240_), .B1(new_n241_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n213_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G230gat), .A2(G233gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT69), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  AOI211_X1 g052(.A(new_n252_), .B(new_n253_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n246_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  OR3_X1    g054(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT68), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(KEYINPUT68), .A3(new_n245_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(new_n253_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT5), .B(G176gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G204gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G120gat), .B(G148gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT70), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n255_), .A2(new_n266_), .A3(new_n258_), .A4(new_n263_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n263_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n202_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  AOI211_X1 g070(.A(KEYINPUT13), .B(new_n269_), .C1(new_n265_), .C2(new_n267_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT103), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G43gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT80), .ZN(new_n276_));
  AND2_X1   g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n278_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT25), .B(G183gat), .ZN(new_n283_));
  INV_X1    g082(.A(G190gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT77), .B1(new_n284_), .B2(KEYINPUT26), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT26), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT26), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(G190gat), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .A4(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT24), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT78), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n290_), .A2(new_n305_), .A3(new_n294_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n301_), .B(new_n302_), .C1(G183gat), .C2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  INV_X1    g111(.A(G176gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(new_n293_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n310_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n307_), .A2(new_n308_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n308_), .B1(new_n307_), .B2(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n282_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n290_), .A2(new_n305_), .A3(new_n294_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n305_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n303_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n317_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT30), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n307_), .A2(new_n308_), .A3(new_n317_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT81), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n281_), .B1(new_n320_), .B2(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n318_), .A2(new_n319_), .A3(new_n282_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n278_), .B(new_n279_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT82), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT81), .B1(new_n325_), .B2(new_n326_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n330_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n281_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT31), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n332_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT82), .B(new_n343_), .C1(new_n328_), .C2(new_n331_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT91), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G204gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G197gat), .ZN(new_n354_));
  INV_X1    g153(.A(G197gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT21), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(G211gat), .A2(G218gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G211gat), .A2(G218gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(KEYINPUT84), .A3(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(KEYINPUT85), .A3(new_n360_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT85), .ZN(new_n364_));
  AND2_X1   g163(.A1(G211gat), .A2(G218gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G211gat), .A2(G218gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n357_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n358_), .A2(new_n371_), .A3(new_n361_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n288_), .A2(G190gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n377_), .A2(new_n286_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n377_), .B2(new_n286_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n283_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n293_), .A2(KEYINPUT24), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(new_n291_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n303_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n314_), .A2(new_n309_), .A3(new_n293_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n376_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n370_), .A2(new_n391_), .A3(new_n374_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n323_), .A2(new_n324_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n375_), .A2(KEYINPUT86), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(new_n307_), .A3(new_n317_), .A4(new_n392_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n389_), .B1(new_n376_), .B2(new_n387_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n352_), .B(new_n399_), .C1(new_n398_), .C2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT97), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT25), .B(G183gat), .Z(new_n408_));
  NOR2_X1   g207(.A1(new_n284_), .A2(KEYINPUT26), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n288_), .A2(G190gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT89), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n377_), .A2(new_n286_), .A3(new_n378_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n294_), .A2(new_n301_), .A3(new_n302_), .A4(new_n298_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n407_), .B(new_n386_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n375_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n407_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT20), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT98), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(KEYINPUT20), .C1(new_n416_), .C2(new_n417_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n395_), .A3(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n422_), .A2(KEYINPUT99), .A3(new_n397_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT99), .B1(new_n422_), .B2(new_n397_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n401_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT100), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n406_), .B1(new_n427_), .B2(new_n352_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n429_));
  INV_X1    g228(.A(G141gat), .ZN(new_n430_));
  INV_X1    g229(.A(G148gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT2), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G155gat), .A2(G162gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n431_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(KEYINPUT1), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n440_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n439_), .A2(KEYINPUT1), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n442_), .B(new_n433_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT29), .ZN(new_n448_));
  XOR2_X1   g247(.A(G22gat), .B(G50gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT28), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n448_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(KEYINPUT29), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n453_));
  OAI211_X1 g252(.A(G228gat), .B(G233gat), .C1(new_n375_), .C2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G78gat), .B(G106gat), .Z(new_n455_));
  NAND2_X1  g254(.A1(G228gat), .A2(G233gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(KEYINPUT83), .A3(KEYINPUT29), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n456_), .B(new_n457_), .C1(new_n393_), .C2(new_n394_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n447_), .B2(KEYINPUT29), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n454_), .B(new_n455_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n451_), .B1(new_n461_), .B2(KEYINPUT88), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n454_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n465_), .A2(KEYINPUT88), .A3(new_n460_), .A4(new_n451_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n403_), .A2(new_n398_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n399_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n351_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT27), .B1(new_n472_), .B2(new_n404_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n345_), .A2(new_n428_), .A3(new_n469_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n340_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n441_), .A2(new_n446_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n340_), .A2(new_n477_), .A3(new_n446_), .A4(new_n441_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(KEYINPUT4), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT4), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n476_), .A2(new_n447_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n482_), .A3(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G57gat), .B(G85gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(G1gat), .B(G29gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n486_), .A2(new_n487_), .A3(new_n493_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT101), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT101), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n488_), .A2(new_n498_), .A3(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n274_), .B1(new_n475_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n422_), .A2(new_n397_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT99), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n422_), .A2(KEYINPUT99), .A3(new_n397_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT100), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n425_), .B(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n405_), .B1(new_n509_), .B2(new_n351_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n342_), .A2(new_n344_), .ZN(new_n511_));
  NOR3_X1   g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n473_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n512_), .A2(KEYINPUT103), .A3(new_n500_), .A4(new_n469_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n502_), .A2(new_n513_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n467_), .A2(new_n468_), .B1(new_n499_), .B2(new_n497_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n428_), .A2(new_n474_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT102), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n351_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n470_), .A2(new_n471_), .A3(new_n519_), .ZN(new_n520_));
  AOI211_X1 g319(.A(new_n500_), .B(new_n520_), .C1(new_n509_), .C2(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n479_), .A2(new_n483_), .A3(new_n480_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n494_), .A2(KEYINPUT95), .A3(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n494_), .A2(new_n522_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT95), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n481_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT96), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  AND4_X1   g328(.A1(new_n523_), .A2(new_n525_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n496_), .A2(KEYINPUT94), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT33), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n472_), .A2(new_n404_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n469_), .B1(new_n521_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n509_), .A2(new_n351_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n473_), .B1(new_n536_), .B2(new_n406_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT102), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n515_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n517_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n511_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n514_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G36gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT73), .B(G29gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT15), .Z(new_n547_));
  XOR2_X1   g346(.A(G1gat), .B(G8gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT74), .ZN(new_n549_));
  INV_X1    g348(.A(G15gat), .ZN(new_n550_));
  INV_X1    g349(.A(G22gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G15gat), .A2(G22gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G1gat), .A2(G8gat), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n552_), .A2(new_n553_), .B1(KEYINPUT14), .B2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n549_), .B(new_n555_), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n546_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n556_), .B(new_n546_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(G229gat), .A3(G233gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT76), .B(G113gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G141gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n561_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n542_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT104), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n542_), .A2(KEYINPUT104), .A3(new_n572_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n273_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n547_), .B2(new_n239_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n546_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n248_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n580_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT72), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n589_), .A3(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  INV_X1    g397(.A(new_n596_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n594_), .A2(new_n595_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n590_), .B(new_n588_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n598_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n213_), .B(new_n607_), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(new_n556_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT16), .B(G183gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(KEYINPUT17), .B2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n609_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n606_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n577_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(G1gat), .A3(new_n500_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n273_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n597_), .A2(new_n601_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n620_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n542_), .A2(new_n572_), .A3(new_n627_), .A4(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n500_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n631_), .ZN(G1324gat));
  OAI21_X1  g431(.A(G8gat), .B1(new_n630_), .B2(new_n537_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(G8gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n537_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n622_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT106), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT106), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT40), .B(new_n634_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  NAND3_X1  g443(.A1(new_n622_), .A2(new_n550_), .A3(new_n345_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G15gat), .B1(new_n630_), .B2(new_n511_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT41), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1326gat));
  OAI21_X1  g447(.A(G22gat), .B1(new_n630_), .B2(new_n469_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n469_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n551_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n623_), .B2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n605_), .A2(KEYINPUT43), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n540_), .A2(new_n511_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n502_), .A2(new_n513_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n604_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(KEYINPUT109), .A3(new_n602_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n514_), .B2(new_n541_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n658_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n572_), .B(new_n620_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT110), .B1(new_n666_), .B2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT44), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT110), .B(new_n672_), .C1(new_n666_), .C2(new_n669_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n500_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n628_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n619_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT104), .B1(new_n542_), .B2(new_n572_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n572_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n574_), .B(new_n679_), .C1(new_n514_), .C2(new_n541_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n627_), .B(new_n677_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n681_), .A2(G29gat), .A3(new_n500_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n675_), .A2(new_n682_), .ZN(G1328gat));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n681_), .A2(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n636_), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n681_), .A2(KEYINPUT111), .A3(G36gat), .A4(new_n537_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n636_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G36gat), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n577_), .A2(new_n692_), .A3(new_n636_), .A4(new_n677_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT111), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n686_), .A2(new_n685_), .A3(new_n636_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(KEYINPUT45), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n689_), .A2(new_n691_), .A3(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n689_), .A2(new_n691_), .A3(new_n696_), .A4(new_n698_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  NOR3_X1   g501(.A1(new_n681_), .A2(G43gat), .A3(new_n511_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n345_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(G43gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g505(.A(G50gat), .B1(new_n674_), .B2(new_n469_), .ZN(new_n707_));
  OR3_X1    g506(.A1(new_n681_), .A2(G50gat), .A3(new_n469_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1331gat));
  NAND2_X1  g508(.A1(new_n273_), .A2(new_n679_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n541_), .B2(new_n514_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n629_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n712_), .A2(G57gat), .A3(new_n501_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n621_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n500_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n713_), .B1(G57gat), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT113), .Z(G1332gat));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n712_), .B2(new_n636_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  INV_X1    g519(.A(new_n714_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n718_), .A3(new_n636_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1333gat));
  NAND2_X1  g522(.A1(new_n712_), .A2(new_n345_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G71gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT114), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT49), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n721_), .A2(new_n345_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n728_), .B(new_n729_), .C1(G71gat), .C2(new_n730_), .ZN(G1334gat));
  INV_X1    g530(.A(G78gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n712_), .B2(new_n652_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT50), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n721_), .A2(new_n732_), .A3(new_n652_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1335gat));
  NOR2_X1   g535(.A1(new_n710_), .A2(new_n619_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n666_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(G85gat), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(new_n500_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n711_), .A2(new_n677_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n501_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n738_), .B2(new_n537_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n636_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(G92gat), .B2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT115), .Z(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n738_), .B2(new_n511_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n741_), .A2(new_n345_), .A3(new_n228_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1338gat));
  OAI21_X1  g551(.A(KEYINPUT117), .B1(new_n738_), .B2(new_n469_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n666_), .A2(new_n754_), .A3(new_n737_), .A4(new_n652_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n757_), .A2(G106gat), .A3(new_n760_), .A4(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n741_), .A2(new_n229_), .A3(new_n652_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n758_), .B(new_n759_), .C1(new_n756_), .C2(new_n229_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n762_), .A2(new_n767_), .A3(new_n764_), .A4(new_n763_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n255_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n246_), .A2(new_n249_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n253_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n246_), .B(KEYINPUT55), .C1(new_n251_), .C2(new_n254_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n262_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n262_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT121), .B(KEYINPUT56), .C1(new_n775_), .C2(new_n262_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n562_), .A2(new_n560_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n559_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n569_), .B(new_n783_), .C1(new_n784_), .C2(new_n560_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(new_n571_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n268_), .A2(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n782_), .A2(KEYINPUT58), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT58), .B1(new_n782_), .B2(new_n787_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n605_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n776_), .A2(KEYINPUT120), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n778_), .A2(new_n779_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n775_), .A2(new_n793_), .A3(KEYINPUT56), .A4(new_n262_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n572_), .A3(new_n268_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n268_), .A2(new_n270_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n786_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n676_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(new_n628_), .C1(new_n796_), .C2(new_n798_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n790_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n679_), .B(new_n619_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT119), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(new_n605_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n804_), .A3(new_n605_), .ZN(new_n808_));
  OAI22_X1  g607(.A1(new_n803_), .A2(new_n619_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n475_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n501_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n572_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(KEYINPUT59), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n809_), .A2(new_n815_), .A3(new_n501_), .A4(new_n810_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n814_), .A2(new_n572_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n817_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g617(.A(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n627_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n812_), .B(new_n820_), .C1(KEYINPUT60), .C2(new_n819_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n814_), .A2(new_n273_), .A3(new_n816_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n819_), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n812_), .B2(new_n619_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n814_), .A2(new_n816_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n619_), .A2(G127gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT122), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1342gat));
  AOI21_X1  g627(.A(G134gat), .B1(new_n812_), .B2(new_n628_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n606_), .A2(G134gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n825_), .B2(new_n830_), .ZN(G1343gat));
  NOR2_X1   g630(.A1(new_n636_), .A2(new_n469_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n809_), .A2(new_n501_), .A3(new_n511_), .A4(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n679_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n430_), .ZN(G1344gat));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n627_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT123), .B(G148gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1345gat));
  NOR2_X1   g637(.A1(new_n833_), .A2(new_n620_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n839_), .B(new_n841_), .ZN(G1346gat));
  INV_X1    g641(.A(new_n833_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G162gat), .B1(new_n843_), .B2(new_n628_), .ZN(new_n844_));
  INV_X1    g643(.A(G162gat), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n663_), .A2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT124), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n843_), .B2(new_n847_), .ZN(G1347gat));
  NOR3_X1   g647(.A1(new_n537_), .A2(new_n501_), .A3(new_n511_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n809_), .A2(new_n469_), .A3(new_n572_), .A4(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G169gat), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n854_));
  INV_X1    g653(.A(new_n312_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n853_), .B(new_n854_), .C1(new_n855_), .C2(new_n850_), .ZN(G1348gat));
  AND2_X1   g655(.A1(new_n809_), .A2(new_n469_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n273_), .A3(new_n849_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n849_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G183gat), .B1(new_n860_), .B2(new_n620_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n619_), .A3(new_n849_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n408_), .B2(new_n862_), .ZN(G1350gat));
  NAND4_X1  g662(.A1(new_n809_), .A2(new_n469_), .A3(new_n606_), .A4(new_n849_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(new_n865_), .A3(G190gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n864_), .B2(G190gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n628_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n860_), .B2(new_n868_), .ZN(G1351gat));
  NAND2_X1  g668(.A1(new_n809_), .A2(new_n511_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n537_), .A2(new_n501_), .A3(new_n469_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n572_), .A3(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n273_), .A3(new_n872_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n353_), .A2(KEYINPUT126), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT127), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n875_), .B(new_n877_), .ZN(G1353gat));
  NAND4_X1  g677(.A1(new_n809_), .A2(new_n511_), .A3(new_n619_), .A4(new_n872_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  AND2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n879_), .B2(new_n880_), .ZN(G1354gat));
  AND2_X1   g682(.A1(new_n871_), .A2(new_n872_), .ZN(new_n884_));
  INV_X1    g683(.A(G218gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n605_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n628_), .A3(new_n872_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n884_), .A2(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1355gat));
endmodule


