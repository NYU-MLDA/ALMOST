//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(KEYINPUT1), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n210_), .B2(KEYINPUT82), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G155gat), .B2(G162gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(new_n207_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n206_), .B1(new_n211_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  INV_X1    g016(.A(G141gat), .ZN(new_n218_));
  INV_X1    g017(.A(G148gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .A4(KEYINPUT83), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n221_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n202_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  INV_X1    g026(.A(new_n207_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n227_), .B1(new_n228_), .B2(new_n209_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n209_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT84), .A3(new_n207_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT85), .B1(new_n216_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT85), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n213_), .A2(new_n214_), .A3(new_n207_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n214_), .B1(new_n213_), .B2(new_n207_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n208_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n234_), .B(new_n235_), .C1(new_n238_), .C2(new_n206_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT29), .B1(new_n233_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G22gat), .B(G50gat), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n241_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n243_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n240_), .A2(new_n241_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n240_), .A2(new_n241_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT29), .B1(new_n216_), .B2(new_n232_), .ZN(new_n250_));
  OR2_X1    g049(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(G204gat), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT90), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT90), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n251_), .A2(new_n256_), .A3(G204gat), .A4(new_n252_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258_));
  INV_X1    g057(.A(G197gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(G204gat), .ZN(new_n260_));
  INV_X1    g059(.A(G204gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n254_), .A2(new_n255_), .A3(new_n257_), .A4(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G211gat), .B(G218gat), .Z(new_n265_));
  NAND3_X1  g064(.A1(new_n251_), .A2(new_n261_), .A3(new_n252_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n255_), .B1(G197gat), .B2(G204gat), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n254_), .A2(new_n257_), .A3(new_n263_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n265_), .A2(KEYINPUT21), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT92), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n264_), .A2(new_n268_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT92), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n250_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G228gat), .A2(G233gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n233_), .A2(KEYINPUT29), .A3(new_n239_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT91), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n269_), .A2(new_n285_), .A3(new_n272_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n233_), .A2(new_n239_), .A3(KEYINPUT87), .A4(KEYINPUT29), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n284_), .A2(new_n288_), .A3(new_n279_), .A4(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G78gat), .B(G106gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n281_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n245_), .B(new_n249_), .C1(new_n294_), .C2(KEYINPUT93), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n281_), .B2(new_n290_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n294_), .A2(new_n296_), .A3(KEYINPUT94), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT94), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n281_), .A2(new_n290_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n291_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n300_), .B2(new_n293_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n295_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT94), .B1(new_n294_), .B2(new_n296_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n249_), .A2(new_n245_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT93), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n293_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n298_), .A3(new_n293_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n303_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n302_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT80), .B(G169gat), .Z(new_n312_));
  NOR2_X1   g111(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT79), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT79), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(G183gat), .A3(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AOI211_X1 g120(.A(new_n315_), .B(new_n316_), .C1(new_n321_), .C2(KEYINPUT23), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT25), .B(G183gat), .ZN(new_n323_));
  INV_X1    g122(.A(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT26), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G190gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(KEYINPUT24), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  INV_X1    g131(.A(G176gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT24), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n328_), .B(new_n331_), .C1(new_n329_), .C2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(G183gat), .B2(G190gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n321_), .B2(new_n336_), .ZN(new_n338_));
  OAI22_X1  g137(.A1(new_n314_), .A2(new_n322_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n273_), .A2(KEYINPUT91), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n275_), .A2(new_n285_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n325_), .A2(new_n327_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT95), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT95), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n323_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n334_), .A2(KEYINPUT96), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT96), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(KEYINPUT24), .C1(new_n332_), .C2(new_n333_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n330_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n316_), .B1(new_n321_), .B2(KEYINPUT23), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n347_), .A2(new_n351_), .A3(new_n352_), .A4(new_n331_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n332_), .A2(new_n333_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G169gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n333_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(new_n338_), .B2(new_n315_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT20), .B1(new_n358_), .B2(new_n275_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n311_), .B1(new_n342_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n340_), .A2(new_n341_), .A3(new_n339_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n311_), .B1(new_n358_), .B2(new_n275_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT20), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n342_), .A2(new_n359_), .A3(new_n311_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n275_), .B(new_n276_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n353_), .A2(new_n357_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT20), .B(new_n361_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n372_), .B2(new_n311_), .ZN(new_n373_));
  OAI211_X1 g172(.A(KEYINPUT27), .B(new_n368_), .C1(new_n373_), .C2(new_n367_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n367_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n361_), .A2(KEYINPUT20), .A3(new_n362_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n311_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n339_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n273_), .B2(new_n371_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n377_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n375_), .B1(new_n376_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n368_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n374_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G71gat), .B(G99gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT81), .B(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n339_), .B(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G127gat), .B(G134gat), .Z(new_n392_));
  XOR2_X1   g191(.A(G113gat), .B(G120gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n391_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT30), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n395_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402_));
  INV_X1    g201(.A(new_n394_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n233_), .A2(new_n239_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n405_), .B(KEYINPUT98), .Z(new_n406_));
  AND2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n233_), .A2(new_n239_), .A3(new_n403_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT97), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n210_), .A2(KEYINPUT82), .ZN(new_n410_));
  INV_X1    g209(.A(new_n208_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n215_), .A3(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n231_), .A2(new_n229_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n412_), .A2(new_n205_), .B1(new_n413_), .B2(new_n226_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n414_), .B2(new_n394_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n205_), .ZN(new_n416_));
  AND4_X1   g215(.A1(new_n409_), .A2(new_n416_), .A3(new_n394_), .A4(new_n235_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n408_), .B(KEYINPUT4), .C1(new_n415_), .C2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n407_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n406_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n408_), .B(new_n420_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT100), .ZN(new_n423_));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n419_), .A2(new_n421_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n401_), .A2(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n309_), .A2(new_n387_), .A3(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n374_), .A2(new_n386_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n303_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n306_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n433_), .B(new_n430_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n418_), .A2(new_n420_), .A3(new_n404_), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n425_), .B(new_n426_), .Z(new_n438_));
  OAI211_X1 g237(.A(new_n408_), .B(new_n406_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n383_), .A2(new_n440_), .A3(new_n368_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n419_), .A2(new_n421_), .A3(new_n427_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT33), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n419_), .A2(new_n444_), .A3(new_n421_), .A4(new_n427_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n441_), .A2(new_n446_), .A3(KEYINPUT101), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT101), .B1(new_n441_), .B2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n360_), .A2(new_n363_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n373_), .A2(new_n449_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n447_), .A2(new_n448_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n436_), .B1(new_n454_), .B2(new_n309_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n401_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n432_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458_));
  INV_X1    g257(.A(G1gat), .ZN(new_n459_));
  INV_X1    g258(.A(G8gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G1gat), .B(G8gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n465_), .A2(KEYINPUT73), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(KEYINPUT73), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n464_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT15), .ZN(new_n477_));
  INV_X1    g276(.A(new_n472_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n469_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(KEYINPUT15), .A3(new_n472_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n464_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n471_), .A2(new_n472_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n464_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n475_), .B1(new_n486_), .B2(new_n473_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G113gat), .B(G141gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT75), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT76), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT77), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n483_), .A2(new_n487_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n491_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT77), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(KEYINPUT76), .A3(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n496_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n492_), .A2(KEYINPUT76), .A3(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(new_n492_), .B2(KEYINPUT76), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n504_), .B(KEYINPUT78), .Z(new_n505_));
  NOR2_X1   g304(.A1(new_n457_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n507_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT10), .B(G99gat), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT9), .ZN(new_n514_));
  INV_X1    g313(.A(G85gat), .ZN(new_n515_));
  INV_X1    g314(.A(G92gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT9), .A3(new_n513_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n510_), .A2(new_n512_), .A3(new_n514_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n513_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT7), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n521_), .B1(KEYINPUT66), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n521_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n520_), .B1(new_n510_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n520_), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT8), .B1(new_n528_), .B2(KEYINPUT67), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n519_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n507_), .B(new_n508_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n528_), .B1(new_n532_), .B2(new_n525_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(new_n529_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n484_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G232gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT34), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n539_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT72), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n542_), .B2(KEYINPUT74), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n480_), .A2(new_n481_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n536_), .B(new_n543_), .C1(new_n544_), .C2(new_n535_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(KEYINPUT74), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n546_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT36), .Z(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n551_), .A2(KEYINPUT36), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n553_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT37), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n464_), .B(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT68), .B(G71gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G78gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n568_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G78gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n567_), .B(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n570_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n566_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n579_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n578_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n564_), .A2(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n512_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n533_), .A2(new_n529_), .B1(new_n590_), .B2(new_n510_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n527_), .A2(new_n530_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n577_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT12), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT64), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n573_), .A2(new_n576_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n531_), .A2(new_n534_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n531_), .B2(new_n534_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(KEYINPUT69), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n595_), .A2(new_n598_), .A3(new_n601_), .A4(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT70), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(KEYINPUT69), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n600_), .B1(new_n608_), .B2(KEYINPUT12), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n609_), .A2(KEYINPUT70), .A3(new_n598_), .A4(new_n604_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n597_), .B1(new_n600_), .B2(new_n593_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n607_), .A2(new_n610_), .A3(new_n611_), .A4(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(KEYINPUT13), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n589_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n506_), .A2(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n626_), .A2(G1gat), .A3(new_n430_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(KEYINPUT104), .B2(KEYINPUT38), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n629_));
  NOR2_X1   g428(.A1(new_n457_), .A2(new_n558_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  INV_X1    g430(.A(new_n504_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n624_), .B2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n622_), .A2(KEYINPUT102), .A3(new_n504_), .A4(new_n623_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(new_n588_), .A3(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n630_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n430_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n638_), .A2(KEYINPUT103), .A3(G1gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT103), .B1(new_n638_), .B2(G1gat), .ZN(new_n640_));
  OAI221_X1 g439(.A(new_n628_), .B1(new_n627_), .B2(new_n629_), .C1(new_n639_), .C2(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n626_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n460_), .A3(new_n387_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n630_), .A2(new_n635_), .A3(new_n645_), .A4(new_n387_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(G8gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n630_), .A2(new_n635_), .A3(new_n387_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT105), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n644_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  AND4_X1   g449(.A1(new_n644_), .A2(new_n649_), .A3(new_n646_), .A4(G8gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n643_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT40), .B(new_n643_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  NAND3_X1  g455(.A1(new_n642_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n636_), .A2(new_n401_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT41), .B1(new_n658_), .B2(G15gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n642_), .A2(new_n662_), .A3(new_n309_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n636_), .A2(new_n309_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(G22gat), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT42), .B(new_n662_), .C1(new_n636_), .C2(new_n309_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n663_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT106), .ZN(G1327gat));
  INV_X1    g468(.A(new_n588_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n558_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n624_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n506_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n637_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n633_), .A2(new_n670_), .A3(new_n634_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n560_), .A2(new_n563_), .A3(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n457_), .A2(new_n680_), .A3(new_n564_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(KEYINPUT43), .ZN(new_n682_));
  INV_X1    g481(.A(new_n432_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n309_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n441_), .A2(new_n446_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n453_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n441_), .A2(new_n446_), .A3(KEYINPUT101), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n387_), .B1(new_n302_), .B2(new_n308_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n684_), .A2(new_n690_), .B1(new_n691_), .B2(new_n430_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n683_), .B1(new_n692_), .B2(new_n401_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n564_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n682_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n677_), .B1(new_n681_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(KEYINPUT108), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n680_), .B1(new_n457_), .B2(new_n564_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n684_), .A2(new_n690_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n401_), .B1(new_n701_), .B2(new_n436_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n694_), .B(new_n682_), .C1(new_n702_), .C2(new_n432_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n676_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n699_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n698_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(KEYINPUT44), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n637_), .A2(G29gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n675_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n433_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n706_), .B2(new_n713_), .ZN(new_n714_));
  AND4_X1   g513(.A1(new_n712_), .A2(new_n506_), .A3(new_n387_), .A4(new_n672_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n716_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n707_), .A2(new_n387_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n705_), .B2(new_n698_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT46), .B(new_n718_), .C1(new_n720_), .C2(new_n712_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n721_), .ZN(G1329gat));
  INV_X1    g521(.A(G43gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n456_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT108), .B1(new_n696_), .B2(new_n697_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n704_), .A2(new_n699_), .A3(KEYINPUT44), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n707_), .B(new_n724_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n673_), .B2(new_n456_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n674_), .B2(new_n309_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n309_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n708_), .B2(new_n734_), .ZN(G1331gat));
  AND2_X1   g534(.A1(new_n622_), .A2(new_n623_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n589_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT110), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n457_), .A2(new_n504_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n637_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n630_), .A2(new_n588_), .A3(new_n624_), .A4(new_n505_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n637_), .B2(KEYINPUT111), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(KEYINPUT111), .B2(new_n743_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n741_), .B1(new_n742_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n742_), .B2(new_n387_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT48), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n740_), .A2(new_n747_), .A3(new_n387_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n740_), .A2(new_n752_), .A3(new_n401_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n742_), .A2(new_n401_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G71gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT49), .B(new_n752_), .C1(new_n742_), .C2(new_n401_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT112), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n753_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1334gat));
  AOI21_X1  g561(.A(new_n574_), .B1(new_n742_), .B2(new_n309_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT50), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n740_), .A2(new_n574_), .A3(new_n309_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1335gat));
  NOR4_X1   g565(.A1(new_n457_), .A2(new_n504_), .A3(new_n736_), .A4(new_n671_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n515_), .A3(new_n637_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n736_), .A2(new_n588_), .A3(new_n504_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(new_n637_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n772_), .B2(new_n515_), .ZN(G1336gat));
  NAND3_X1  g572(.A1(new_n767_), .A2(new_n516_), .A3(new_n387_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n771_), .A2(new_n387_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n516_), .ZN(G1337gat));
  INV_X1    g575(.A(new_n511_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n401_), .A3(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n771_), .A2(new_n401_), .ZN(new_n779_));
  INV_X1    g578(.A(G99gat), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT113), .B(new_n778_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g581(.A(G106gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n767_), .A2(new_n783_), .A3(new_n309_), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT52), .B(new_n783_), .C1(new_n771_), .C2(new_n309_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n309_), .B(new_n769_), .C1(new_n681_), .C2(new_n695_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g589(.A(G113gat), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n505_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n736_), .A2(new_n505_), .A3(new_n564_), .A4(new_n588_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT115), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n794_), .B(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(new_n473_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n482_), .A2(new_n800_), .A3(new_n475_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n486_), .A2(new_n473_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n801_), .B(new_n496_), .C1(new_n802_), .C2(new_n475_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n492_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n799_), .B1(new_n620_), .B2(new_n805_), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT118), .B(new_n804_), .C1(new_n617_), .C2(new_n619_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n504_), .A2(new_n619_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT116), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n504_), .A2(new_n619_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n605_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n598_), .B1(new_n609_), .B2(new_n604_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n607_), .A2(new_n610_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n616_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n618_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n810_), .B(new_n812_), .C1(new_n820_), .C2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n808_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n562_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n820_), .A2(new_n822_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n619_), .A2(new_n805_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n564_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(KEYINPUT57), .A3(new_n562_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n827_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n798_), .B1(new_n838_), .B2(new_n670_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n684_), .A2(new_n637_), .A3(new_n433_), .A4(new_n401_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT120), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n793_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n824_), .B2(new_n562_), .ZN(new_n844_));
  AOI211_X1 g643(.A(new_n826_), .B(new_n558_), .C1(new_n808_), .C2(new_n823_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n588_), .B1(new_n846_), .B2(new_n836_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT59), .B(new_n841_), .C1(new_n847_), .C2(new_n798_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n792_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n839_), .A2(new_n632_), .A3(new_n842_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n850_), .A2(new_n851_), .A3(G113gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n850_), .B2(G113gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n852_), .B2(new_n853_), .ZN(G1340gat));
  NOR2_X1   g653(.A1(new_n839_), .A2(new_n842_), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n736_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n855_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n856_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n736_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n856_), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n861_), .A3(new_n588_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n670_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1342gat));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n855_), .A2(new_n865_), .A3(new_n558_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n564_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1343gat));
  NAND3_X1  g667(.A1(new_n691_), .A2(new_n637_), .A3(new_n456_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n839_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n504_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n624_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g673(.A1(new_n870_), .A2(new_n588_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  NOR3_X1   g676(.A1(new_n839_), .A2(new_n562_), .A3(new_n869_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT122), .B1(new_n878_), .B2(G162gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n564_), .A2(new_n881_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n882_), .A2(new_n883_), .B1(new_n870_), .B2(new_n884_), .ZN(G1347gat));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n309_), .A2(new_n433_), .A3(new_n431_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n839_), .A2(new_n632_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n886_), .B1(new_n889_), .B2(new_n332_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n504_), .B(new_n887_), .C1(new_n847_), .C2(new_n798_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(KEYINPUT62), .A3(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n355_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n891_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT123), .B1(new_n891_), .B2(G169gat), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n893_), .A2(new_n898_), .ZN(G1348gat));
  NOR2_X1   g698(.A1(new_n839_), .A2(new_n888_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n624_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n588_), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n323_), .B(G183gat), .S(new_n903_), .Z(G1350gat));
  NAND4_X1  g703(.A1(new_n900_), .A2(new_n345_), .A3(new_n346_), .A4(new_n558_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n839_), .A2(new_n564_), .A3(new_n888_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n324_), .ZN(G1351gat));
  NAND3_X1  g706(.A1(new_n309_), .A2(new_n430_), .A3(new_n456_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n908_), .A2(KEYINPUT124), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(KEYINPUT124), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n433_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n839_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n504_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n624_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT125), .B(G204gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1353gat));
  NOR3_X1   g717(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n913_), .A2(new_n588_), .A3(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(KEYINPUT127), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n921_), .B(new_n923_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n913_), .A2(new_n925_), .A3(new_n558_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n839_), .A2(new_n564_), .A3(new_n912_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n925_), .ZN(G1355gat));
endmodule


