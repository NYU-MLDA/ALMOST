//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209_));
  OAI211_X1 g008(.A(KEYINPUT21), .B(new_n207_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  INV_X1    g010(.A(new_n208_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(KEYINPUT92), .ZN(new_n213_));
  XOR2_X1   g012(.A(G197gat), .B(G204gat), .Z(new_n214_));
  OAI21_X1  g013(.A(new_n214_), .B1(KEYINPUT21), .B2(new_n208_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n210_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT81), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT22), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n219_), .A2(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT82), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G176gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n217_), .B1(new_n223_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT83), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(new_n217_), .C1(new_n223_), .C2(new_n229_), .ZN(new_n233_));
  INV_X1    g032(.A(G183gat), .ZN(new_n234_));
  INV_X1    g033(.A(G190gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT23), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(G183gat), .A3(G190gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(KEYINPUT84), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT84), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n240_), .B(KEYINPUT23), .C1(new_n234_), .C2(new_n235_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n239_), .B(new_n241_), .C1(G183gat), .C2(G190gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n231_), .A2(new_n233_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244_));
  NAND2_X1  g043(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT26), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n234_), .A2(KEYINPUT25), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G183gat), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .A4(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT80), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT80), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n252_), .A2(new_n258_), .A3(new_n255_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT24), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n236_), .A2(new_n238_), .B1(new_n260_), .B2(new_n253_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n243_), .A2(new_n244_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n244_), .B1(new_n243_), .B2(new_n262_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n216_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n253_), .A2(new_n260_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n239_), .A2(new_n269_), .A3(new_n241_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT95), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n239_), .A2(KEYINPUT95), .A3(new_n269_), .A4(new_n241_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n249_), .A2(new_n251_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n247_), .A2(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n235_), .A2(KEYINPUT26), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT94), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n274_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n272_), .A2(new_n255_), .A3(new_n273_), .A4(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n216_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n217_), .B(KEYINPUT96), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n226_), .A2(new_n228_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n224_), .A2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n236_), .A2(new_n238_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  OAI221_X1 g087(.A(new_n283_), .B1(new_n284_), .B2(new_n286_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n290_), .A2(KEYINPUT20), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n265_), .A2(new_n268_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n243_), .A2(new_n262_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT85), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n243_), .A2(new_n244_), .A3(new_n262_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n282_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n281_), .A2(new_n289_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n297_), .B1(new_n298_), .B2(new_n216_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n268_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n206_), .B1(new_n292_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT97), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n263_), .A2(new_n264_), .A3(new_n216_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n216_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT20), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n267_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n265_), .A2(new_n291_), .A3(new_n268_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n205_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n302_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT97), .B(new_n206_), .C1(new_n292_), .C2(new_n300_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT100), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(KEYINPUT100), .A3(new_n310_), .A4(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n303_), .A2(new_n305_), .A3(new_n267_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n268_), .B1(new_n265_), .B2(new_n291_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n206_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT27), .A3(new_n308_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G57gat), .B(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT98), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G155gat), .B(G162gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT90), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT2), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(KEYINPUT90), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G141gat), .ZN(new_n337_));
  INV_X1    g136(.A(G148gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT3), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n334_), .A2(new_n336_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342_));
  AND4_X1   g141(.A1(KEYINPUT89), .A2(new_n342_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT89), .B1(new_n344_), .B2(new_n342_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n331_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n339_), .A2(new_n348_), .A3(new_n332_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(KEYINPUT1), .B2(new_n330_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  INV_X1    g151(.A(G134gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G127gat), .ZN(new_n354_));
  INV_X1    g153(.A(G127gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G134gat), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT86), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT86), .B1(new_n354_), .B2(new_n356_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G113gat), .B(G120gat), .Z(new_n361_));
  INV_X1    g160(.A(KEYINPUT86), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n355_), .A2(G134gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n353_), .A2(G127gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT86), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n361_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n352_), .B1(new_n360_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT87), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n351_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n347_), .B(new_n350_), .C1(new_n360_), .C2(new_n367_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n371_), .A2(KEYINPUT4), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n351_), .A2(new_n368_), .A3(new_n370_), .A4(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n329_), .B1(new_n373_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n371_), .A2(KEYINPUT4), .A3(new_n372_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(KEYINPUT98), .A3(new_n377_), .A4(new_n375_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n328_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n379_), .A2(new_n327_), .A3(new_n383_), .A4(new_n382_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n282_), .B1(KEYINPUT29), .B2(new_n351_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G228gat), .A2(G233gat), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G78gat), .B(G106gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n351_), .A2(KEYINPUT29), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n400_));
  XNOR2_X1  g199(.A(G22gat), .B(G50gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n399_), .B(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n396_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(KEYINPUT93), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n395_), .A2(new_n397_), .A3(KEYINPUT93), .A4(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410_));
  INV_X1    g209(.A(G43gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT31), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n263_), .A2(new_n264_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(G15gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT30), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n368_), .A2(new_n370_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n415_), .A2(new_n419_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n414_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n423_), .A3(new_n413_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n322_), .A2(new_n388_), .A3(new_n409_), .A4(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT101), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n408_), .A2(new_n320_), .A3(new_n388_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n316_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n309_), .A2(new_n311_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n382_), .A2(new_n383_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT33), .A3(new_n327_), .A4(new_n379_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n386_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n381_), .A2(new_n376_), .A3(new_n375_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n371_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n328_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n438_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n306_), .A2(new_n307_), .A3(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n317_), .A2(new_n318_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n387_), .B(new_n447_), .C1(new_n448_), .C2(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n409_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n435_), .A2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT88), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT88), .B1(new_n426_), .B2(new_n428_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n432_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n433_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n408_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n455_), .B(new_n432_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n431_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G29gat), .B(G36gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT72), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT72), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n463_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471_));
  INV_X1    g270(.A(G1gat), .ZN(new_n472_));
  INV_X1    g271(.A(G8gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G1gat), .B(G8gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n470_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT77), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n470_), .B(KEYINPUT15), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n477_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n470_), .A2(new_n478_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n481_), .B(KEYINPUT78), .Z(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G141gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  AND3_X1   g290(.A1(new_n483_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G85gat), .B(G92gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT67), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT8), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT6), .Z(new_n500_));
  NOR2_X1   g299(.A1(G99gat), .A2(G106gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT7), .Z(new_n502_));
  OAI21_X1  g301(.A(new_n496_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n500_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n495_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT10), .B(G99gat), .Z(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT65), .B(G85gat), .Z(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(new_n506_), .A3(G92gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n505_), .A2(new_n507_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n498_), .A2(new_n503_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n504_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n484_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n504_), .A2(new_n470_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G232gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT34), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT73), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n517_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n520_), .A2(new_n521_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT36), .Z(new_n535_));
  AND2_X1   g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(new_n537_), .A3(new_n530_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT37), .B1(new_n536_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n535_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT37), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n538_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT11), .ZN(new_n547_));
  XOR2_X1   g346(.A(G71gat), .B(G78gat), .Z(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n546_), .A2(KEYINPUT11), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n548_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT68), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n515_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT64), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT68), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n552_), .B(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n561_), .A2(new_n504_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n549_), .B(KEYINPUT12), .C1(new_n550_), .C2(new_n551_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n515_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n557_), .A2(new_n559_), .A3(new_n562_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n554_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n559_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n578_), .B1(new_n581_), .B2(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n477_), .B(new_n585_), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n552_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT75), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G183gat), .B(G211gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(KEYINPUT17), .A3(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT76), .Z(new_n595_));
  XOR2_X1   g394(.A(new_n593_), .B(KEYINPUT17), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n586_), .B(new_n553_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n545_), .A2(new_n584_), .A3(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n461_), .A2(new_n494_), .A3(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT102), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n472_), .A3(new_n387_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n461_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n536_), .A2(new_n539_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n583_), .A2(new_n494_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n599_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT103), .Z(new_n611_));
  AND2_X1   g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n388_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n603_), .A2(new_n604_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n605_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n602_), .A2(new_n473_), .A3(new_n321_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n612_), .A2(new_n321_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n618_), .A2(G8gat), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n618_), .B2(G8gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(G1325gat));
  INV_X1    g423(.A(new_n455_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n417_), .B1(new_n612_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT41), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n417_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n601_), .B2(new_n628_), .ZN(G1326gat));
  OAI21_X1  g428(.A(G22gat), .B1(new_n613_), .B2(new_n409_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n409_), .A2(G22gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n601_), .B2(new_n632_), .ZN(G1327gat));
  INV_X1    g432(.A(new_n494_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n607_), .A2(new_n599_), .ZN(new_n635_));
  NOR4_X1   g434(.A1(new_n606_), .A2(new_n634_), .A3(new_n584_), .A4(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n387_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n599_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n609_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n544_), .B(KEYINPUT105), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n461_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n545_), .A2(new_n641_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n459_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n644_), .B1(new_n647_), .B2(new_n431_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n640_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT44), .B(new_n640_), .C1(new_n643_), .C2(new_n648_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n387_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT106), .B1(new_n656_), .B2(G29gat), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n638_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(G36gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n636_), .A2(new_n660_), .A3(new_n321_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT45), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n651_), .A2(new_n321_), .A3(new_n653_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n663_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT107), .B1(new_n663_), .B2(G36gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n662_), .B(new_n667_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  NOR4_X1   g470(.A1(new_n652_), .A2(new_n654_), .A3(new_n411_), .A4(new_n429_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G43gat), .B1(new_n636_), .B2(new_n625_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n672_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n636_), .B2(new_n408_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n408_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n655_), .B2(new_n680_), .ZN(G1331gat));
  NOR2_X1   g480(.A1(new_n606_), .A2(new_n494_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n682_), .A2(new_n584_), .A3(new_n639_), .A4(new_n544_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT110), .ZN(new_n684_));
  AOI21_X1  g483(.A(G57gat), .B1(new_n684_), .B2(new_n387_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n583_), .A2(new_n494_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n608_), .A2(new_n639_), .A3(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT111), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n387_), .B2(KEYINPUT112), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(KEYINPUT112), .B2(new_n689_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n688_), .B2(new_n691_), .ZN(G1332gat));
  INV_X1    g491(.A(G64gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n693_), .A3(new_n321_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n688_), .A2(new_n321_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(G64gat), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT48), .B(new_n693_), .C1(new_n688_), .C2(new_n321_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  NOR2_X1   g498(.A1(new_n455_), .A2(G71gat), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT114), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n684_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n688_), .A2(new_n625_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(G71gat), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G71gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n684_), .A2(new_n708_), .A3(new_n408_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT50), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n688_), .A2(new_n408_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G78gat), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT50), .B(new_n708_), .C1(new_n688_), .C2(new_n408_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1335gat));
  NAND4_X1  g513(.A1(new_n682_), .A2(new_n584_), .A3(new_n599_), .A4(new_n607_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n387_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n686_), .A2(new_n599_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n643_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n648_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT115), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n387_), .A2(new_n511_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(G1336gat));
  INV_X1    g523(.A(G92gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n716_), .A2(new_n725_), .A3(new_n321_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n722_), .A2(new_n321_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n725_), .ZN(G1337gat));
  NAND2_X1  g527(.A1(new_n721_), .A2(new_n625_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G99gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n716_), .A2(new_n430_), .A3(new_n508_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n716_), .A2(new_n509_), .A3(new_n408_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n721_), .A2(new_n408_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G106gat), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT52), .B(new_n509_), .C1(new_n721_), .C2(new_n408_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g540(.A(KEYINPUT118), .ZN(new_n742_));
  INV_X1    g541(.A(new_n574_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n562_), .A2(new_n565_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n555_), .B1(new_n515_), .B2(new_n553_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n568_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n566_), .B2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n744_), .A2(new_n745_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT55), .B1(new_n749_), .B2(new_n559_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n743_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT56), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n485_), .A2(new_n486_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(KEYINPUT117), .ZN(new_n754_));
  INV_X1    g553(.A(new_n487_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(KEYINPUT117), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n491_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n492_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n743_), .C1(new_n748_), .C2(new_n750_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n752_), .A2(new_n759_), .A3(new_n575_), .A4(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT58), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n576_), .B1(new_n751_), .B2(KEYINPUT56), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n759_), .A4(new_n761_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n742_), .B1(new_n767_), .B2(new_n545_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n494_), .A3(new_n761_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n759_), .A2(new_n578_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n607_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT57), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n607_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n768_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n767_), .A2(new_n545_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT118), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n639_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n583_), .A2(new_n544_), .A3(new_n634_), .A4(new_n639_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT54), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT119), .B1(new_n780_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n768_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n773_), .A2(new_n775_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n599_), .B1(new_n787_), .B2(new_n778_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n782_), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n321_), .A2(new_n388_), .A3(new_n408_), .A4(new_n429_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n784_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(G113gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n494_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n786_), .A2(new_n777_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n783_), .B1(new_n599_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n792_), .B2(KEYINPUT59), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(new_n494_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n795_), .B1(new_n802_), .B2(new_n794_), .ZN(G1340gat));
  INV_X1    g602(.A(G120gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n801_), .B2(new_n584_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n583_), .B2(KEYINPUT60), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(KEYINPUT60), .B2(new_n804_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n792_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT120), .B1(new_n805_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810_));
  INV_X1    g609(.A(new_n808_), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n583_), .B(new_n800_), .C1(new_n792_), .C2(KEYINPUT59), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n810_), .B(new_n811_), .C1(new_n812_), .C2(new_n804_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n793_), .B2(new_n639_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n355_), .B1(new_n639_), .B2(KEYINPUT121), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(KEYINPUT121), .B2(new_n355_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n815_), .B1(new_n801_), .B2(new_n817_), .ZN(G1342gat));
  NAND3_X1  g617(.A1(new_n793_), .A2(new_n353_), .A3(new_n607_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n801_), .A2(new_n545_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n353_), .ZN(G1343gat));
  AND2_X1   g620(.A1(new_n784_), .A2(new_n790_), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n625_), .A2(new_n321_), .A3(new_n388_), .A4(new_n409_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n634_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(new_n337_), .ZN(G1344gat));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n583_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT122), .B(G148gat), .Z(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(G1345gat));
  NOR2_X1   g628(.A1(new_n824_), .A2(new_n599_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT61), .B(G155gat), .Z(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1346gat));
  INV_X1    g631(.A(new_n824_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n833_), .A2(G162gat), .A3(new_n642_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G162gat), .B1(new_n833_), .B2(new_n607_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1347gat));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n322_), .A2(new_n387_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n625_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n408_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n797_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n494_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n837_), .B1(new_n843_), .B2(G169gat), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT62), .B(new_n221_), .C1(new_n842_), .C2(new_n494_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n797_), .A2(KEYINPUT123), .A3(new_n841_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n494_), .A2(new_n224_), .A3(new_n285_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n844_), .A2(new_n845_), .B1(new_n849_), .B2(new_n850_), .ZN(G1348gat));
  INV_X1    g650(.A(new_n284_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n584_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n822_), .A2(new_n409_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n839_), .A2(new_n225_), .A3(new_n583_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n852_), .A2(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(G1349gat));
  NOR3_X1   g655(.A1(new_n849_), .A2(new_n274_), .A3(new_n599_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n854_), .A2(new_n625_), .A3(new_n639_), .A4(new_n838_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n234_), .ZN(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n849_), .B2(new_n544_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n607_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT124), .Z(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n849_), .B2(new_n862_), .ZN(G1351gat));
  NOR4_X1   g662(.A1(new_n322_), .A2(new_n625_), .A3(new_n387_), .A4(new_n409_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n784_), .A2(new_n790_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n494_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n584_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT63), .B(G211gat), .Z(new_n871_));
  NAND4_X1  g670(.A1(new_n865_), .A2(new_n870_), .A3(new_n639_), .A4(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n784_), .A2(new_n790_), .A3(new_n639_), .A4(new_n864_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n871_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT125), .B1(new_n873_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n872_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n872_), .A2(new_n877_), .A3(KEYINPUT126), .A4(new_n875_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1354gat));
  NAND2_X1  g681(.A1(new_n865_), .A2(new_n607_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT127), .B(G218gat), .Z(new_n884_));
  NOR2_X1   g683(.A1(new_n544_), .A2(new_n884_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(new_n865_), .B2(new_n885_), .ZN(G1355gat));
endmodule


