//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_;
  XNOR2_X1  g000(.A(KEYINPUT88), .B(G204gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G197gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G197gat), .B2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206_));
  NOR3_X1   g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n202_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT89), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G197gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n213_), .A2(G204gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n211_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n205_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n204_), .A2(KEYINPUT90), .A3(new_n205_), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT90), .B1(new_n204_), .B2(new_n205_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n206_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n208_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT24), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT96), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT96), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT24), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT95), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n239_), .A2(new_n232_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n235_), .A2(new_n236_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n228_), .A2(new_n224_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(G183gat), .B2(G190gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G169gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n231_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n237_), .A3(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n222_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n229_), .B1(G183gat), .B2(G190gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT22), .B1(new_n254_), .B2(new_n230_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n231_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n237_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT78), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(new_n259_), .B2(G183gat), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n260_), .B(new_n241_), .C1(new_n240_), .C2(new_n258_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n232_), .A2(KEYINPUT24), .A3(new_n237_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n244_), .A4(new_n233_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n221_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n250_), .A2(KEYINPUT20), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT93), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n264_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n279_), .B(new_n208_), .C1(new_n217_), .C2(new_n220_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n280_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n222_), .A2(new_n249_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT94), .B1(new_n280_), .B2(KEYINPUT20), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n272_), .B(new_n278_), .C1(new_n284_), .C2(new_n270_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT82), .Z(new_n287_));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  OR2_X1    g088(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n289_), .A2(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT84), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n287_), .B(new_n288_), .C1(new_n296_), .C2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n288_), .B(KEYINPUT1), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n287_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G113gat), .B(G120gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n299_), .A2(new_n302_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT85), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n305_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n308_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(KEYINPUT4), .A3(new_n313_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n315_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n310_), .B(new_n304_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n308_), .A2(KEYINPUT4), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT0), .ZN(new_n325_));
  INV_X1    g124(.A(G57gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n323_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n316_), .A2(new_n322_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n285_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n266_), .A2(new_n270_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n284_), .B2(new_n271_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT98), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n278_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n284_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n336_), .B1(new_n341_), .B2(new_n270_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT98), .B1(new_n342_), .B2(new_n277_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n335_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT99), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT99), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n335_), .B(new_n346_), .C1(new_n340_), .C2(new_n343_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(KEYINPUT97), .A3(new_n276_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n314_), .A2(new_n318_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n317_), .A2(new_n315_), .A3(new_n321_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n329_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n332_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n352_), .B2(new_n332_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT97), .ZN(new_n355_));
  INV_X1    g154(.A(new_n276_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n338_), .B2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n338_), .A2(new_n356_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n348_), .B(new_n354_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n345_), .A2(new_n347_), .A3(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n305_), .A2(new_n311_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n363_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n364_), .B1(new_n363_), .B2(new_n367_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT87), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n303_), .A2(new_n366_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n222_), .B2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n221_), .B(new_n374_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n372_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n381_), .A3(new_n371_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n370_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n386_), .A3(new_n370_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n264_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393_));
  INV_X1    g192(.A(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n395_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n392_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n392_), .A2(new_n400_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n308_), .B(KEYINPUT31), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT81), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n390_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n272_), .B1(new_n270_), .B2(new_n284_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(new_n276_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n358_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n348_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n414_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n333_), .A2(KEYINPUT100), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n333_), .A2(KEYINPUT100), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n388_), .A2(new_n410_), .A3(new_n389_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n408_), .A2(new_n409_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n389_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n387_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n420_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n360_), .A2(new_n411_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G230gat), .A2(G233gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G99gat), .A2(G106gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT6), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT10), .B(G99gat), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT64), .B(G92gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT9), .B1(new_n434_), .B2(G85gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  OAI221_X1 g237(.A(new_n430_), .B1(G106gat), .B2(new_n432_), .C1(new_n435_), .C2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G85gat), .B(G92gat), .ZN(new_n441_));
  INV_X1    g240(.A(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(G106gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT67), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT66), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT7), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT66), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT67), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT66), .B(new_n446_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  AOI211_X1 g253(.A(KEYINPUT8), .B(new_n441_), .C1(new_n454_), .C2(new_n430_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n450_), .A2(KEYINPUT68), .A3(new_n453_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT68), .B1(new_n450_), .B2(new_n453_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n430_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n441_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n456_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT69), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n455_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n430_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT68), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n448_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT7), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n448_), .B1(new_n447_), .B2(KEYINPUT67), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AOI211_X1 g268(.A(KEYINPUT7), .B(new_n448_), .C1(new_n447_), .C2(KEYINPUT67), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n465_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n450_), .A2(KEYINPUT68), .A3(new_n453_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n464_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT8), .B1(new_n473_), .B2(new_n441_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT69), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n440_), .B1(new_n463_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G57gat), .B(G64gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n478_));
  XOR2_X1   g277(.A(G71gat), .B(G78gat), .Z(new_n479_));
  NOR2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n479_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n477_), .A2(KEYINPUT11), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n428_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n462_), .B(KEYINPUT8), .C1(new_n473_), .C2(new_n441_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n455_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n459_), .A2(new_n460_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n462_), .B1(new_n489_), .B2(KEYINPUT8), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n439_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n492_));
  INV_X1    g291(.A(new_n484_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n485_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n439_), .B(new_n484_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT70), .B1(new_n476_), .B2(new_n484_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n500_), .A3(new_n493_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n498_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n496_), .B1(new_n502_), .B2(new_n427_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G120gat), .B(G148gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT5), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G176gat), .B(G204gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n507_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n496_), .B(new_n509_), .C1(new_n502_), .C2(new_n427_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT13), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n515_), .A2(KEYINPUT71), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(KEYINPUT71), .ZN(new_n517_));
  XOR2_X1   g316(.A(G43gat), .B(G50gat), .Z(new_n518_));
  OR3_X1    g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT15), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(KEYINPUT15), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G8gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n522_), .A2(new_n523_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT77), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n521_), .A2(new_n530_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT76), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n522_), .A2(KEYINPUT77), .A3(new_n523_), .A4(new_n530_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n521_), .A2(new_n530_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n535_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n543_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n514_), .A2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n522_), .A2(new_n523_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n491_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT72), .ZN(new_n553_));
  INV_X1    g352(.A(new_n521_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT34), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n476_), .A2(new_n554_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT72), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n491_), .A2(new_n560_), .A3(new_n551_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n553_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n558_), .A2(new_n555_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT36), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n553_), .A2(new_n559_), .A3(new_n569_), .A4(new_n561_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT73), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT73), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n564_), .A2(new_n573_), .A3(new_n568_), .A4(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n564_), .A2(new_n570_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n567_), .B(KEYINPUT36), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT75), .ZN(new_n587_));
  XOR2_X1   g386(.A(G183gat), .B(G211gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(KEYINPUT17), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(KEYINPUT17), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n530_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n484_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n591_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n575_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n584_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n426_), .A2(new_n550_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n525_), .A3(new_n420_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT38), .Z(new_n603_));
  INV_X1    g402(.A(new_n579_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n339_), .B1(new_n338_), .B2(new_n278_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n342_), .A2(KEYINPUT98), .A3(new_n277_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n334_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n359_), .B1(new_n607_), .B2(new_n346_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n347_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n411_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n417_), .A2(new_n425_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n604_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n550_), .A2(new_n597_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n525_), .B1(new_n614_), .B2(new_n420_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n603_), .A2(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n417_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n601_), .A2(new_n526_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n612_), .A2(new_n619_), .A3(new_n617_), .A4(new_n613_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(G8gat), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n617_), .A3(new_n613_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT101), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n621_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n622_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n618_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(KEYINPUT40), .B(new_n618_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1325gat));
  AOI21_X1  g430(.A(new_n397_), .B1(new_n614_), .B2(new_n410_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n601_), .A2(new_n397_), .A3(new_n410_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n614_), .B2(new_n390_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT42), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n601_), .A2(new_n638_), .A3(new_n390_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  AND2_X1   g441(.A1(new_n584_), .A2(new_n599_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT43), .B1(new_n426_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n610_), .A2(new_n611_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n643_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n514_), .A2(new_n549_), .A3(new_n597_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(G29gat), .A3(new_n420_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n644_), .B2(new_n648_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT44), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n426_), .A2(new_n550_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n579_), .A2(new_n598_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n419_), .B2(new_n418_), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n653_), .A2(new_n655_), .B1(G29gat), .B2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT102), .ZN(G1328gat));
  NAND2_X1  g460(.A1(new_n652_), .A2(new_n617_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G36gat), .B1(new_n662_), .B2(new_n655_), .ZN(new_n663_));
  INV_X1    g462(.A(G36gat), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n656_), .A2(new_n664_), .A3(new_n617_), .A4(new_n657_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n663_), .A2(new_n666_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1329gat));
  OAI21_X1  g470(.A(new_n394_), .B1(new_n658_), .B2(new_n422_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n652_), .A2(G43gat), .A3(new_n410_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(new_n655_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g474(.A(new_n658_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G50gat), .B1(new_n676_), .B2(new_n390_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n652_), .A2(G50gat), .A3(new_n390_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n654_), .A2(KEYINPUT44), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n426_), .A2(new_n549_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT104), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n514_), .B1(new_n681_), .B2(KEYINPUT104), .ZN(new_n683_));
  INV_X1    g482(.A(new_n600_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n420_), .A4(new_n684_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(KEYINPUT105), .A3(new_n326_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT105), .B1(new_n685_), .B2(new_n326_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n514_), .ZN(new_n688_));
  AND4_X1   g487(.A1(new_n612_), .A2(new_n548_), .A3(new_n688_), .A4(new_n598_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT106), .B(G57gat), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n420_), .A3(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n686_), .A2(new_n687_), .A3(new_n691_), .ZN(G1332gat));
  AND2_X1   g491(.A1(new_n682_), .A2(new_n683_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n684_), .ZN(new_n694_));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n617_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n689_), .B2(new_n617_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT48), .Z(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1333gat));
  INV_X1    g498(.A(G71gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n700_), .A3(new_n410_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n689_), .B2(new_n410_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n703_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT107), .B(KEYINPUT49), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n704_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n701_), .B1(new_n707_), .B2(new_n708_), .ZN(G1334gat));
  INV_X1    g508(.A(G78gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n694_), .A2(new_n710_), .A3(new_n390_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n689_), .B2(new_n390_), .ZN(new_n712_));
  XOR2_X1   g511(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1335gat));
  NAND3_X1  g514(.A1(new_n688_), .A2(new_n548_), .A3(new_n597_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT110), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n649_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n420_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G85gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n682_), .A2(new_n657_), .A3(new_n683_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n420_), .A2(new_n328_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(G1336gat));
  NAND3_X1  g522(.A1(new_n693_), .A2(new_n617_), .A3(new_n657_), .ZN(new_n724_));
  INV_X1    g523(.A(G92gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n617_), .A2(new_n434_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT111), .ZN(new_n727_));
  AOI22_X1  g526(.A1(new_n724_), .A2(new_n725_), .B1(new_n718_), .B2(new_n727_), .ZN(G1337gat));
  NOR3_X1   g527(.A1(new_n721_), .A2(new_n432_), .A3(new_n422_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n442_), .B1(new_n718_), .B2(new_n410_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(KEYINPUT112), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n729_), .A2(new_n730_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1338gat));
  NAND3_X1  g534(.A1(new_n649_), .A2(new_n390_), .A3(new_n717_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G106gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n390_), .A2(new_n443_), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n738_), .A2(new_n739_), .B1(new_n721_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  OAI221_X1 g542(.A(new_n743_), .B1(new_n721_), .B2(new_n740_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  AOI21_X1  g544(.A(new_n549_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n643_), .A2(KEYINPUT54), .A3(new_n598_), .A4(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748_));
  INV_X1    g547(.A(new_n746_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n600_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n546_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n537_), .A2(KEYINPUT115), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n537_), .A2(KEYINPUT115), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n540_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n535_), .A2(new_n541_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n547_), .B1(new_n757_), .B2(new_n538_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n476_), .A2(KEYINPUT70), .A3(new_n484_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n500_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n497_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n428_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n509_), .B1(new_n763_), .B2(new_n496_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n510_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n759_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT116), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n511_), .A2(new_n768_), .A3(new_n759_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n497_), .A2(new_n427_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT12), .B1(new_n476_), .B2(new_n484_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n498_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(KEYINPUT55), .A2(new_n774_), .B1(new_n775_), .B2(new_n427_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n496_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT56), .B(new_n507_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n507_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n496_), .A2(new_n777_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n774_), .A2(KEYINPUT55), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n786_), .B(new_n787_), .C1(new_n427_), .C2(new_n775_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n784_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n788_), .A2(new_n781_), .A3(new_n507_), .A4(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n780_), .A2(new_n785_), .A3(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n548_), .A2(new_n765_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n770_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n752_), .B1(new_n793_), .B2(new_n604_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n792_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n767_), .A2(new_n769_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n797_), .A2(KEYINPUT57), .A3(new_n579_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n779_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n507_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n510_), .B(new_n759_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n584_), .A2(new_n599_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n794_), .A2(new_n798_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n751_), .B1(new_n806_), .B2(new_n597_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n417_), .A2(new_n420_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n421_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT117), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n549_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n807_), .B2(new_n810_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n809_), .B(KEYINPUT117), .Z(new_n816_));
  AOI21_X1  g615(.A(new_n604_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n817_), .A2(KEYINPUT57), .B1(new_n803_), .B2(new_n804_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n598_), .B1(new_n818_), .B2(new_n794_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(KEYINPUT59), .C1(new_n819_), .C2(new_n751_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n548_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n813_), .B1(new_n821_), .B2(new_n812_), .ZN(G1340gat));
  AOI21_X1  g621(.A(new_n514_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n823_));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  INV_X1    g623(.A(new_n811_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n514_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n823_), .A2(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1341gat));
  INV_X1    g627(.A(G127gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n811_), .A2(new_n829_), .A3(new_n598_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n597_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n829_), .ZN(G1342gat));
  NAND2_X1  g631(.A1(new_n815_), .A2(new_n820_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n646_), .A2(G134gat), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT118), .Z(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n811_), .A2(new_n604_), .ZN(new_n839_));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n837_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n835_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G134gat), .B1(new_n811_), .B2(new_n604_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT119), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n845_), .ZN(G1343gat));
  NOR2_X1   g645(.A1(new_n808_), .A2(new_n424_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT120), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n807_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n549_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n688_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT121), .B(G148gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1345gat));
  NAND2_X1  g653(.A1(new_n849_), .A2(new_n598_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  NOR2_X1   g656(.A1(new_n579_), .A2(G162gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n849_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G162gat), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n807_), .A2(new_n643_), .A3(new_n848_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n859_), .B(KEYINPUT122), .C1(new_n860_), .C2(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n420_), .A2(new_n422_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n617_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n617_), .B2(new_n868_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n389_), .B(new_n388_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n807_), .A2(new_n548_), .A3(new_n872_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n874_));
  OR3_X1    g673(.A1(new_n873_), .A2(new_n230_), .A3(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n230_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n246_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  NOR2_X1   g677(.A1(new_n807_), .A2(new_n872_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n688_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n598_), .ZN(new_n882_));
  MUX2_X1   g681(.A(new_n240_), .B(G183gat), .S(new_n882_), .Z(G1350gat));
  NAND3_X1  g682(.A1(new_n879_), .A2(new_n604_), .A3(new_n241_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n646_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(new_n886_), .A3(G190gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n885_), .B2(G190gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(G1351gat));
  NOR3_X1   g688(.A1(new_n417_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n807_), .A2(new_n548_), .A3(new_n891_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n892_), .A2(KEYINPUT126), .A3(G197gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(G197gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT126), .B1(new_n892_), .B2(G197gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1352gat));
  NOR2_X1   g695(.A1(new_n807_), .A2(new_n891_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n209_), .A4(new_n688_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n688_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT127), .B1(new_n900_), .B2(G204gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n202_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n899_), .B1(new_n901_), .B2(new_n902_), .ZN(G1353gat));
  INV_X1    g702(.A(new_n897_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n904_), .A2(new_n597_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT63), .B(G211gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n897_), .A2(new_n598_), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1354gat));
  OR3_X1    g707(.A1(new_n904_), .A2(G218gat), .A3(new_n579_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G218gat), .B1(new_n904_), .B2(new_n643_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1355gat));
endmodule


