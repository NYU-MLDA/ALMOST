//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT23), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n207_), .A2(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n208_), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT81), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT25), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n218_), .B(new_n221_), .C1(new_n222_), .C2(new_n219_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n214_), .A2(new_n205_), .A3(KEYINPUT81), .A4(new_n206_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n213_), .A2(new_n217_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(new_n211_), .B2(new_n209_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(new_n211_), .B2(new_n209_), .ZN(new_n228_));
  OAI21_X1  g027(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n225_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT83), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n233_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT31), .ZN(new_n237_));
  XOR2_X1   g036(.A(G71gat), .B(G99gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G15gat), .B(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT82), .B(KEYINPUT30), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n242_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n237_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G197gat), .A2(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G197gat), .A2(G204gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT21), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  AND2_X1   g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(new_n252_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G211gat), .B(G218gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n257_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n225_), .A2(new_n264_), .A3(new_n232_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n222_), .A2(new_n218_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n213_), .A2(new_n215_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n232_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n264_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT90), .B1(new_n265_), .B2(KEYINPUT20), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n251_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n264_), .A2(new_n268_), .A3(new_n232_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT91), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n233_), .A2(new_n270_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n251_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n278_), .A2(KEYINPUT20), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n264_), .A2(new_n268_), .A3(new_n280_), .A4(new_n232_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n276_), .A2(new_n277_), .A3(new_n279_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G8gat), .B(G36gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT18), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n274_), .A2(new_n287_), .A3(new_n282_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  INV_X1    g091(.A(new_n282_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n265_), .A2(KEYINPUT20), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT90), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(new_n271_), .A3(new_n266_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n293_), .B1(new_n297_), .B2(new_n251_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n292_), .B1(new_n298_), .B2(new_n287_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n296_), .A2(new_n278_), .A3(new_n271_), .A4(new_n266_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n277_), .A2(KEYINPUT20), .A3(new_n275_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n251_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n288_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n291_), .A2(new_n292_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT84), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  NOR4_X1   g110(.A1(KEYINPUT85), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT2), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G141gat), .A3(G148gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G141gat), .ZN(new_n323_));
  INV_X1    g122(.A(G148gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT3), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n311_), .B1(new_n317_), .B2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n315_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT85), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n314_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n319_), .A2(new_n321_), .B1(new_n325_), .B2(KEYINPUT3), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT86), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n310_), .B1(new_n328_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n309_), .B(KEYINPUT1), .Z(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n308_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n337_), .A2(new_n325_), .A3(new_n318_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT87), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n310_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n332_), .A2(KEYINPUT86), .A3(new_n333_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT86), .B1(new_n332_), .B2(new_n333_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n337_), .A2(new_n325_), .A3(new_n318_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT29), .B1(new_n339_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G22gat), .B(G50gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT28), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n270_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n357_), .B(KEYINPUT29), .C1(new_n335_), .C2(new_n338_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n339_), .A2(new_n346_), .A3(KEYINPUT29), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n264_), .A2(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n352_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n350_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n364_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT29), .B1(new_n335_), .B2(new_n338_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n264_), .B1(new_n369_), .B2(KEYINPUT88), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n353_), .B1(new_n370_), .B2(new_n359_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n351_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(new_n352_), .A3(new_n364_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n367_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n339_), .A2(new_n346_), .A3(new_n246_), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n245_), .B(KEYINPUT92), .Z(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G1gat), .B(G29gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT93), .B(G85gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT0), .B(G57gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n376_), .A2(KEYINPUT4), .A3(new_n378_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n339_), .A2(new_n346_), .A3(new_n387_), .A4(new_n246_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n379_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n380_), .B(new_n385_), .C1(new_n386_), .C2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n376_), .A2(new_n378_), .A3(KEYINPUT4), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(new_n389_), .A3(new_n388_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n385_), .B1(new_n394_), .B2(new_n380_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n372_), .A2(new_n373_), .A3(new_n366_), .A4(new_n350_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n305_), .A2(new_n375_), .A3(new_n396_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT33), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n391_), .A2(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n274_), .A2(new_n287_), .A3(new_n282_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n287_), .B1(new_n274_), .B2(new_n282_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n394_), .A2(KEYINPUT33), .A3(new_n380_), .A4(new_n385_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n393_), .A2(new_n379_), .A3(new_n388_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n385_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n376_), .A2(new_n378_), .A3(new_n389_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n298_), .B2(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n375_), .A2(new_n397_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n398_), .A2(KEYINPUT94), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n292_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n304_), .A2(KEYINPUT27), .A3(new_n290_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n380_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n406_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n391_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT94), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n397_), .A4(new_n375_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n249_), .B1(new_n416_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n248_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n415_), .A2(new_n305_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G29gat), .B(G36gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT71), .ZN(new_n432_));
  INV_X1    g231(.A(G36gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G29gat), .ZN(new_n434_));
  INV_X1    g233(.A(G29gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G36gat), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n434_), .A2(new_n436_), .A3(KEYINPUT71), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n431_), .A2(KEYINPUT71), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n442_), .B2(new_n437_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n440_), .A2(new_n443_), .A3(KEYINPUT15), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT15), .B1(new_n440_), .B2(new_n443_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447_));
  INV_X1    g246(.A(G1gat), .ZN(new_n448_));
  INV_X1    g247(.A(G8gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G8gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n440_), .A2(new_n443_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G229gat), .A2(G233gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT76), .Z(new_n459_));
  NAND3_X1  g258(.A1(new_n454_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n455_), .B(new_n456_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G229gat), .A3(G233gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G113gat), .B(G141gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT77), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G169gat), .B(G197gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  AND3_X1   g266(.A1(new_n463_), .A2(KEYINPUT78), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n467_), .B1(new_n463_), .B2(KEYINPUT78), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n430_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n472_));
  XOR2_X1   g271(.A(G85gat), .B(G92gat), .Z(new_n473_));
  INV_X1    g272(.A(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT64), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n474_), .A3(new_n475_), .A4(KEYINPUT64), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n473_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT10), .B(G99gat), .Z(new_n487_));
  AOI22_X1  g286(.A1(KEYINPUT9), .A2(new_n473_), .B1(new_n487_), .B2(new_n475_), .ZN(new_n488_));
  INV_X1    g287(.A(G85gat), .ZN(new_n489_));
  INV_X1    g288(.A(G92gat), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT9), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n483_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n473_), .A2(KEYINPUT8), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n480_), .B2(KEYINPUT65), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n477_), .A2(new_n497_), .A3(new_n479_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n472_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n480_), .A2(KEYINPUT65), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n481_), .B(KEYINPUT6), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(KEYINPUT8), .A3(new_n473_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n484_), .A2(new_n485_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT66), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n509_));
  XOR2_X1   g308(.A(G71gat), .B(G78gat), .Z(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n509_), .A2(new_n510_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n500_), .A2(new_n506_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n505_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n515_), .A2(KEYINPUT12), .A3(new_n512_), .A4(new_n511_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n513_), .B1(new_n500_), .B2(new_n506_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n514_), .B(new_n516_), .C1(new_n517_), .C2(KEYINPUT12), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G230gat), .A2(G233gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n514_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n522_), .B2(new_n517_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G120gat), .B(G148gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT5), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n521_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT67), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n521_), .A2(new_n523_), .A3(new_n531_), .A4(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n521_), .A2(new_n523_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n527_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT13), .B1(new_n533_), .B2(new_n535_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n513_), .B(new_n453_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G127gat), .B(G155gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT16), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G183gat), .B(G211gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n545_), .A2(new_n546_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n541_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT75), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT75), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n500_), .A2(new_n456_), .A3(new_n506_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT69), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n446_), .B2(new_n515_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n559_), .A2(new_n563_), .A3(KEYINPUT35), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n559_), .B2(KEYINPUT35), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n446_), .A2(new_n515_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(KEYINPUT72), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT72), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n446_), .B2(new_n515_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n555_), .B(new_n561_), .C1(new_n571_), .C2(new_n566_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT36), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n569_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n575_), .B(KEYINPUT36), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT37), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT73), .B(KEYINPUT37), .C1(new_n577_), .C2(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n569_), .A2(new_n572_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n569_), .A2(KEYINPUT74), .A3(new_n572_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n578_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT37), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n569_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n554_), .B1(new_n585_), .B2(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n471_), .A2(new_n538_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n448_), .A3(new_n422_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  INV_X1    g396(.A(new_n554_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n470_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n538_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n592_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT95), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n601_), .B1(new_n430_), .B2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n417_), .A2(new_n421_), .A3(new_n418_), .A4(new_n391_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT94), .B1(new_n415_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n414_), .A2(new_n415_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n607_), .A2(new_n425_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n248_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n428_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT96), .A3(new_n603_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n600_), .B1(new_n605_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n396_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n597_), .A2(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n595_), .A2(new_n449_), .A3(new_n419_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n419_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(G8gat), .ZN(new_n620_));
  AOI211_X1 g419(.A(KEYINPUT39), .B(new_n449_), .C1(new_n613_), .C2(new_n419_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(G1325gat));
  INV_X1    g423(.A(G15gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n595_), .A2(new_n625_), .A3(new_n249_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G15gat), .B1(new_n614_), .B2(new_n248_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT41), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(G1326gat));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n415_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n595_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n613_), .A2(new_n633_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(G22gat), .ZN(new_n637_));
  AOI211_X1 g436(.A(KEYINPUT42), .B(new_n632_), .C1(new_n613_), .C2(new_n633_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT97), .ZN(G1327gat));
  INV_X1    g439(.A(new_n602_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n554_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT100), .Z(new_n643_));
  OR2_X1    g442(.A1(new_n536_), .A2(new_n537_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n471_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n435_), .A3(new_n422_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n586_), .A2(new_n578_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n592_), .ZN(new_n651_));
  AOI21_X1  g450(.A(KEYINPUT73), .B1(new_n651_), .B2(KEYINPUT37), .ZN(new_n652_));
  INV_X1    g451(.A(new_n584_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT98), .B(new_n593_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT98), .B1(new_n585_), .B2(new_n593_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n585_), .A2(new_n593_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n658_), .A2(KEYINPUT43), .B1(new_n611_), .B2(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n644_), .A2(new_n598_), .A3(new_n470_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n649_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n661_), .B1(new_n611_), .B2(new_n657_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n610_), .B2(new_n428_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n665_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n422_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n672_), .A2(KEYINPUT99), .A3(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT99), .B1(new_n672_), .B2(G29gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n648_), .B1(new_n673_), .B2(new_n674_), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n646_), .A2(G36gat), .A3(new_n305_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n667_), .A2(new_n419_), .A3(new_n670_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT101), .B1(new_n679_), .B2(G36gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  OAI221_X1 g484(.A(new_n678_), .B1(new_n683_), .B2(KEYINPUT46), .C1(new_n680_), .C2(new_n681_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  INV_X1    g486(.A(G43gat), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n248_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n667_), .A2(new_n670_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n667_), .A2(KEYINPUT103), .A3(new_n670_), .A4(new_n689_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n646_), .B2(new_n248_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g495(.A(G50gat), .B1(new_n647_), .B2(new_n633_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n633_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n671_), .B2(new_n698_), .ZN(G1331gat));
  NOR3_X1   g498(.A1(new_n430_), .A2(new_n599_), .A3(new_n538_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n594_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT104), .Z(new_n702_));
  AOI21_X1  g501(.A(G57gat), .B1(new_n702_), .B2(new_n422_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n644_), .A2(new_n598_), .A3(new_n470_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n605_), .B2(new_n612_), .ZN(new_n705_));
  INV_X1    g504(.A(G57gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n422_), .B2(KEYINPUT105), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(KEYINPUT105), .B2(new_n706_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n705_), .B2(new_n708_), .ZN(G1332gat));
  NOR2_X1   g508(.A1(new_n305_), .A2(G64gat), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT106), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n702_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n705_), .A2(new_n419_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G64gat), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n713_), .A3(G64gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n249_), .A2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT107), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n702_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT49), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n705_), .A2(new_n249_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G71gat), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT49), .B(new_n718_), .C1(new_n705_), .C2(new_n249_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n702_), .A2(new_n727_), .A3(new_n633_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n705_), .A2(new_n633_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G78gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT50), .B(new_n727_), .C1(new_n705_), .C2(new_n633_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1335gat));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n598_), .A2(new_n599_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n644_), .B2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n735_), .B(new_n734_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n664_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n396_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n643_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n700_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n489_), .A3(new_n422_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n741_), .B2(new_n305_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n490_), .A3(new_n419_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n741_), .B2(new_n248_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n249_), .A2(new_n487_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n744_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n753_), .B(new_n754_), .Z(G1338gat));
  NAND3_X1  g554(.A1(new_n745_), .A2(new_n475_), .A3(new_n633_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n740_), .A2(new_n633_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G106gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT52), .B(new_n475_), .C1(new_n740_), .C2(new_n633_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g561(.A1(new_n538_), .A2(new_n594_), .A3(new_n470_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT54), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n538_), .A2(new_n594_), .A3(new_n767_), .A4(new_n470_), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n768_), .A2(KEYINPUT110), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n763_), .A2(KEYINPUT111), .A3(KEYINPUT54), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(KEYINPUT110), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n766_), .A2(new_n769_), .A3(new_n770_), .A4(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n533_), .A2(new_n535_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n463_), .A2(new_n467_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n461_), .A2(new_n459_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT113), .B1(new_n775_), .B2(new_n467_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n459_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n454_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(KEYINPUT113), .A3(new_n467_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n774_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n470_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n520_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n519_), .A2(KEYINPUT55), .ZN(new_n785_));
  OR3_X1    g584(.A1(new_n518_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n518_), .A2(new_n784_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n527_), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n786_), .A2(KEYINPUT56), .A3(new_n527_), .A4(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n773_), .A2(new_n780_), .B1(new_n781_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n641_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(new_n641_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n533_), .A3(new_n780_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT58), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n660_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(KEYINPUT58), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n795_), .B(new_n796_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n554_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n772_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n633_), .A2(new_n419_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n422_), .A3(new_n249_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT59), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n809_), .B(new_n806_), .C1(new_n772_), .C2(new_n803_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(G113gat), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n470_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n804_), .A2(new_n807_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n815_), .B2(new_n470_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT115), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n813_), .C1(new_n815_), .C2(new_n470_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n812_), .A2(new_n814_), .B1(new_n817_), .B2(new_n819_), .ZN(G1340gat));
  OAI21_X1  g619(.A(G120gat), .B1(new_n811_), .B2(new_n538_), .ZN(new_n821_));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n538_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(KEYINPUT60), .B2(new_n822_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n821_), .B1(new_n815_), .B2(new_n824_), .ZN(G1341gat));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n815_), .B2(new_n554_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n598_), .A2(G127gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT116), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n826_), .B(new_n828_), .C1(new_n811_), .C2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n763_), .A2(KEYINPUT111), .A3(KEYINPUT54), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT111), .B1(new_n763_), .B2(KEYINPUT54), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n768_), .B(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n835_), .A2(new_n837_), .B1(new_n802_), .B2(new_n554_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n809_), .B1(new_n838_), .B2(new_n806_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n804_), .A2(KEYINPUT59), .A3(new_n807_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n831_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n806_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G127gat), .B1(new_n842_), .B2(new_n598_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT117), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n832_), .A2(new_n844_), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n815_), .B2(new_n603_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n660_), .A2(G134gat), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT118), .B(new_n847_), .C1(new_n811_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G134gat), .B1(new_n842_), .B2(new_n604_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1343gat));
  NAND4_X1  g653(.A1(new_n633_), .A2(new_n422_), .A3(new_n305_), .A4(new_n248_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT119), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n772_), .B2(new_n803_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n599_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT120), .B(G141gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n644_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n598_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n858_), .A2(KEYINPUT121), .A3(new_n598_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n858_), .B2(new_n604_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n657_), .A2(G162gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n858_), .B2(new_n873_), .ZN(G1347gat));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n415_), .A2(new_n419_), .A3(new_n427_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n838_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n599_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n878_), .B2(G169gat), .ZN(new_n879_));
  AOI211_X1 g678(.A(KEYINPUT62), .B(new_n203_), .C1(new_n877_), .C2(new_n599_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n876_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT122), .B1(new_n804_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n883_), .B(new_n876_), .C1(new_n772_), .C2(new_n803_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n230_), .A2(new_n203_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n599_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n879_), .A2(new_n880_), .B1(new_n885_), .B2(new_n888_), .ZN(G1348gat));
  NAND2_X1  g688(.A1(new_n804_), .A2(new_n881_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G176gat), .B1(new_n890_), .B2(new_n538_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n644_), .A2(new_n204_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n885_), .B2(new_n892_), .ZN(G1349gat));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n220_), .B1(new_n890_), .B2(new_n554_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n554_), .A2(new_n222_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n894_), .B(new_n895_), .C1(new_n885_), .C2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n883_), .B1(new_n838_), .B2(new_n876_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n804_), .A2(KEYINPUT122), .A3(new_n881_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G183gat), .B1(new_n877_), .B2(new_n598_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT123), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n898_), .A2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n885_), .B2(new_n659_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n604_), .A2(new_n218_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n885_), .B2(new_n906_), .ZN(G1351gat));
  NAND3_X1  g706(.A1(new_n633_), .A2(new_n396_), .A3(new_n248_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n419_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n909_), .B2(new_n908_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n804_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n599_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n538_), .ZN(new_n916_));
  INV_X1    g715(.A(G204gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(KEYINPUT125), .B2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT125), .B(G204gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n916_), .B2(new_n919_), .ZN(G1353gat));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921_));
  INV_X1    g720(.A(G211gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n598_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT126), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n913_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n922_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1354gat));
  OR3_X1    g726(.A1(new_n912_), .A2(G218gat), .A3(new_n603_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G218gat), .B1(new_n912_), .B2(new_n659_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1355gat));
endmodule


