//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(KEYINPUT7), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT65), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT64), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n209_), .B(new_n204_), .C1(new_n211_), .C2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n205_), .A2(KEYINPUT7), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n206_), .A2(new_n208_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(KEYINPUT10), .B(G99gat), .Z(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT9), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G85gat), .A3(G92gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .A4(new_n208_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n220_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n216_), .A2(new_n217_), .A3(new_n229_), .A4(new_n218_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n221_), .A2(new_n228_), .A3(new_n230_), .A4(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT67), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n221_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n202_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI211_X1 g044(.A(KEYINPUT68), .B(new_n202_), .C1(new_n239_), .C2(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT12), .B1(new_n240_), .B2(new_n241_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n240_), .A2(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n221_), .A2(KEYINPUT69), .A3(new_n228_), .A4(new_n230_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(KEYINPUT12), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n247_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n238_), .A2(new_n202_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT70), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  NOR4_X1   g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n247_), .A4(new_n255_), .ZN(new_n260_));
  OAI22_X1  g059(.A1(new_n245_), .A2(new_n246_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G120gat), .B(G148gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(G204gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT5), .ZN(new_n264_));
  INV_X1    g063(.A(G176gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n257_), .A2(new_n260_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n202_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n238_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n242_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT68), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n243_), .A2(new_n244_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n266_), .B1(new_n269_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT13), .B1(new_n268_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n261_), .A2(new_n267_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n269_), .A2(new_n277_), .A3(new_n266_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G113gat), .B(G141gat), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G197gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(G29gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G15gat), .B(G22gat), .Z(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT77), .B(G8gat), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G1gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n298_), .B2(KEYINPUT14), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT78), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G1gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n299_), .B(KEYINPUT78), .ZN(new_n303_));
  INV_X1    g102(.A(G1gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n302_), .A2(new_n305_), .A3(G8gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(G8gat), .B1(new_n302_), .B2(new_n305_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n295_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n303_), .A2(new_n304_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n301_), .A2(G1gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT15), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n295_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n302_), .A2(new_n305_), .A3(G8gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n308_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n295_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n320_), .A3(new_n316_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n308_), .B2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n291_), .B1(new_n319_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n318_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n306_), .A2(new_n307_), .A3(new_n295_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n308_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n291_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n323_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT16), .B(G183gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G211gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G155gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT17), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n306_), .A2(new_n307_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G231gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n237_), .B(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n337_), .B1(new_n343_), .B2(KEYINPUT79), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345_));
  INV_X1    g144(.A(new_n337_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n341_), .A2(new_n345_), .A3(new_n342_), .A4(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n336_), .A2(KEYINPUT17), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n344_), .A2(new_n347_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G190gat), .B(G218gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G134gat), .ZN(new_n352_));
  INV_X1    g151(.A(G162gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(KEYINPUT36), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G232gat), .A2(G233gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT72), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT34), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT75), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n363_), .A2(KEYINPUT75), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n314_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n362_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n240_), .B2(new_n320_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n364_), .B(new_n365_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n251_), .A2(new_n315_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n368_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT75), .A4(new_n363_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n357_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n369_), .A2(new_n372_), .A3(new_n357_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n374_), .A2(new_n375_), .B1(KEYINPUT36), .B2(new_n355_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT37), .B1(new_n373_), .B2(KEYINPUT76), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n355_), .A2(KEYINPUT36), .ZN(new_n380_));
  INV_X1    g179(.A(new_n375_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n373_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(new_n377_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n350_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G197gat), .A2(G204gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT91), .B(G204gat), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT21), .B(new_n385_), .C1(new_n386_), .C2(G197gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(G211gat), .B(G218gat), .Z(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n290_), .A2(G204gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n386_), .B2(new_n290_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n387_), .B(new_n389_), .C1(new_n391_), .C2(KEYINPUT21), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT21), .A3(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT26), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT26), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n401_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G183gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT25), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(G183gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT80), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n400_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n288_), .A2(new_n265_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  NOR2_X1   g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT82), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(new_n410_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n414_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421_));
  INV_X1    g220(.A(G190gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n404_), .B2(new_n422_), .ZN(new_n423_));
  AND4_X1   g222(.A1(new_n414_), .A2(new_n423_), .A3(new_n419_), .A4(new_n415_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  OR3_X1    g224(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT25), .B(G183gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n402_), .B1(new_n428_), .B2(KEYINPUT80), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n426_), .B(new_n427_), .C1(new_n429_), .C2(new_n400_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n413_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n418_), .B1(G183gat), .B2(G190gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n409_), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT22), .B(G169gat), .Z(new_n434_));
  OAI211_X1 g233(.A(new_n432_), .B(new_n433_), .C1(G176gat), .C2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n395_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT26), .B(G190gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n412_), .B1(new_n438_), .B2(new_n428_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n435_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n394_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n436_), .A2(KEYINPUT20), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT19), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n441_), .A2(new_n394_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n431_), .A2(new_n435_), .ZN(new_n449_));
  AOI211_X1 g248(.A(new_n447_), .B(new_n448_), .C1(new_n449_), .C2(new_n394_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n450_), .B2(new_n445_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G8gat), .B(G36gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  AND2_X1   g255(.A1(new_n451_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT96), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT27), .ZN(new_n459_));
  INV_X1    g258(.A(new_n445_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n443_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n450_), .B2(new_n460_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n456_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n451_), .A2(new_n456_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT96), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G155gat), .B(G162gat), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(KEYINPUT1), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471_));
  INV_X1    g270(.A(G141gat), .ZN(new_n472_));
  INV_X1    g271(.A(G148gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G141gat), .A2(G148gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(new_n470_), .A2(new_n471_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n471_), .B1(new_n470_), .B2(new_n477_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n469_), .B(KEYINPUT88), .Z(new_n481_));
  OR2_X1    g280(.A1(new_n474_), .A2(KEYINPUT3), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT2), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(KEYINPUT3), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n480_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G127gat), .B(G134gat), .ZN(new_n490_));
  INV_X1    g289(.A(G113gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G120gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n478_), .A2(new_n479_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n495_));
  INV_X1    g294(.A(G120gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n492_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n498_), .A3(KEYINPUT93), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(KEYINPUT4), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n494_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT94), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n499_), .A2(new_n501_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n506_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT0), .B(G57gat), .ZN(new_n511_));
  INV_X1    g310(.A(G85gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G1gat), .B(G29gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n505_), .A2(new_n507_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(new_n516_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n451_), .A2(new_n456_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n459_), .B1(new_n457_), .B2(new_n522_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n468_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G227gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT84), .ZN(new_n527_));
  INV_X1    g326(.A(G71gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G99gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT30), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n431_), .A2(new_n532_), .A3(new_n435_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G15gat), .B(G43gat), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n449_), .A2(KEYINPUT30), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n431_), .A2(new_n532_), .A3(new_n435_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n531_), .B1(new_n536_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n535_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n530_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n525_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(new_n525_), .A3(new_n544_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n493_), .B(KEYINPUT31), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n546_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n542_), .A2(new_n543_), .A3(new_n530_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n530_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT85), .ZN(new_n555_));
  INV_X1    g354(.A(new_n549_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT86), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n545_), .A3(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G22gat), .B(G50gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT28), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(KEYINPUT90), .A2(G233gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(G228gat), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT29), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n495_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n569_), .B2(new_n395_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n394_), .B(new_n566_), .C1(new_n495_), .C2(new_n568_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT89), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n489_), .A2(KEYINPUT29), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G78gat), .B(G106gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  AOI21_X1  g376(.A(new_n572_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n574_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n575_), .B(new_n576_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n578_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n573_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n562_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n577_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(new_n580_), .A3(new_n573_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n561_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n552_), .A2(new_n559_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n552_), .B2(new_n559_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n524_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n457_), .A2(new_n522_), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n517_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n519_), .B(new_n516_), .C1(new_n594_), .C2(KEYINPUT33), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n505_), .A2(new_n506_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n516_), .B1(new_n509_), .B2(new_n507_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n591_), .A2(new_n593_), .A3(new_n595_), .A4(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT32), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n451_), .B1(new_n600_), .B2(new_n463_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n462_), .A2(KEYINPUT32), .A3(new_n456_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n601_), .B(new_n602_), .C1(new_n518_), .C2(new_n520_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n559_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n552_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n604_), .B(new_n587_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n384_), .B1(new_n590_), .B2(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n286_), .A2(new_n331_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n521_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n304_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT97), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616_));
  INV_X1    g415(.A(new_n283_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n282_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n331_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT98), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n284_), .A2(new_n621_), .A3(new_n331_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n616_), .B1(new_n624_), .B2(new_n349_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n382_), .B(KEYINPUT100), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n590_), .B2(new_n607_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(KEYINPUT99), .A3(new_n350_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n521_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n614_), .A2(new_n615_), .A3(new_n630_), .ZN(G1324gat));
  NAND2_X1  g430(.A1(new_n468_), .A2(new_n523_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n297_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n609_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n625_), .A2(new_n632_), .A3(new_n627_), .A4(new_n628_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT39), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(G8gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n635_), .B2(G8gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g439(.A(G15gat), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n606_), .A2(new_n605_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n609_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n629_), .A2(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(new_n645_), .B2(G15gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(G1326gat));
  XNOR2_X1  g447(.A(new_n587_), .B(KEYINPUT101), .ZN(new_n649_));
  OAI21_X1  g448(.A(G22gat), .B1(new_n629_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT103), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n653_), .ZN(new_n655_));
  INV_X1    g454(.A(G22gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n649_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n609_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(new_n655_), .A3(new_n658_), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n350_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n590_), .A2(new_n607_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n376_), .A2(new_n378_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n382_), .A2(new_n377_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n661_), .B1(new_n662_), .B2(new_n666_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT43), .B(new_n665_), .C1(new_n590_), .C2(new_n607_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n660_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n660_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n521_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n662_), .A2(new_n626_), .A3(new_n349_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(new_n331_), .A3(new_n284_), .ZN(new_n678_));
  INV_X1    g477(.A(G29gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n610_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(G36gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n682_), .A3(new_n632_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n675_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n682_), .B1(new_n686_), .B2(new_n632_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT46), .ZN(G1329gat));
  OAI21_X1  g488(.A(G43gat), .B1(new_n675_), .B2(new_n644_), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n678_), .A2(new_n691_), .A3(new_n642_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g493(.A(new_n587_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n672_), .A2(new_n695_), .A3(new_n674_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n672_), .A2(KEYINPUT106), .A3(new_n695_), .A4(new_n674_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(G50gat), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n698_), .A2(KEYINPUT107), .A3(G50gat), .A4(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(G50gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n678_), .A2(new_n705_), .A3(new_n657_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(KEYINPUT108), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1331gat));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n331_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n608_), .A2(new_n713_), .A3(new_n279_), .A4(new_n283_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT109), .Z(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n716_), .B2(new_n521_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n286_), .A2(new_n331_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n627_), .A3(new_n350_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT110), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(KEYINPUT111), .B2(G57gat), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n712_), .B1(new_n610_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT112), .Z(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n715_), .A2(new_n726_), .A3(new_n632_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n632_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G64gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT48), .B(new_n726_), .C1(new_n720_), .C2(new_n632_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  NAND3_X1  g531(.A1(new_n715_), .A2(new_n528_), .A3(new_n642_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n720_), .A2(new_n642_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G71gat), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT49), .B(new_n528_), .C1(new_n720_), .C2(new_n642_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  INV_X1    g537(.A(G78gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n715_), .A2(new_n739_), .A3(new_n657_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n720_), .A2(new_n657_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G78gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT50), .B(new_n739_), .C1(new_n720_), .C2(new_n657_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n718_), .A2(new_n677_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n610_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n667_), .A2(new_n668_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n749_), .A2(new_n331_), .A3(new_n284_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n349_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n521_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n752_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n747_), .B2(new_n632_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n632_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(G92gat), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n747_), .A2(new_n222_), .A3(new_n642_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G99gat), .B1(new_n751_), .B2(new_n644_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n759_), .A2(new_n760_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n758_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n747_), .A2(new_n223_), .A3(new_n695_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  INV_X1    g568(.A(new_n751_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n695_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(G106gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT52), .B(new_n223_), .C1(new_n770_), .C2(new_n695_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n768_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  AND3_X1   g577(.A1(new_n254_), .A2(KEYINPUT117), .A3(new_n239_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT117), .B1(new_n254_), .B2(new_n239_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n270_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n254_), .A2(KEYINPUT55), .A3(new_n256_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n267_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n318_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n308_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n291_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n330_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n268_), .A2(new_n795_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n785_), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(new_n267_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n791_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n665_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n791_), .A2(new_n798_), .A3(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n791_), .A2(new_n798_), .A3(new_n804_), .A4(KEYINPUT58), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n801_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n268_), .A2(new_n278_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(new_n795_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n281_), .A2(new_n331_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n788_), .A2(new_n790_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  OAI22_X1  g614(.A1(new_n813_), .A2(new_n626_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n815_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n809_), .B(KEYINPUT116), .ZN(new_n818_));
  INV_X1    g617(.A(new_n790_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n267_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n818_), .A2(new_n821_), .B1(new_n807_), .B2(new_n795_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n626_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n822_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n806_), .A2(new_n816_), .A3(new_n817_), .A4(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n349_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n331_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n349_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT115), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n837_), .B(new_n834_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n830_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n713_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n840_), .B2(new_n384_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n837_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n833_), .A2(KEYINPUT115), .A3(new_n835_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n829_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n826_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n632_), .A2(new_n521_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n588_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n845_), .B1(new_n825_), .B2(new_n349_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT121), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n849_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n331_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n853_), .A2(new_n851_), .A3(new_n858_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n713_), .B(new_n859_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g660(.A(new_n496_), .B1(new_n284_), .B2(KEYINPUT60), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n856_), .B(new_n862_), .C1(KEYINPUT60), .C2(new_n496_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n286_), .B(new_n859_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n496_), .ZN(G1341gat));
  AOI21_X1  g664(.A(G127gat), .B1(new_n856_), .B2(new_n350_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n859_), .B1(new_n855_), .B2(KEYINPUT59), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n350_), .A2(G127gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT123), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n867_), .B2(new_n869_), .ZN(G1342gat));
  AOI21_X1  g669(.A(G134gat), .B1(new_n856_), .B2(new_n626_), .ZN(new_n871_));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n872_), .B(new_n859_), .C1(new_n855_), .C2(KEYINPUT59), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n666_), .ZN(G1343gat));
  AND3_X1   g673(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n846_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT121), .B1(new_n826_), .B2(new_n846_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n589_), .A3(new_n850_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G141gat), .B1(new_n878_), .B2(new_n713_), .ZN(new_n879_));
  AND4_X1   g678(.A1(new_n589_), .A2(new_n849_), .A3(new_n850_), .A4(new_n854_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n472_), .A3(new_n331_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1344gat));
  OAI21_X1  g681(.A(G148gat), .B1(new_n878_), .B2(new_n286_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n286_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n473_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1345gat));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT124), .Z(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n878_), .B2(new_n349_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n880_), .A2(new_n350_), .A3(new_n888_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1346gat));
  NOR3_X1   g691(.A1(new_n878_), .A2(new_n353_), .A3(new_n665_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G162gat), .B1(new_n880_), .B2(new_n626_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n847_), .A2(new_n649_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n755_), .A2(new_n610_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n642_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n713_), .A2(new_n434_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT125), .Z(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n331_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(G169gat), .ZN(new_n905_));
  AOI211_X1 g704(.A(KEYINPUT62), .B(new_n288_), .C1(new_n899_), .C2(new_n331_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n902_), .B1(new_n905_), .B2(new_n906_), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n877_), .A2(new_n587_), .A3(new_n884_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G176gat), .B1(new_n908_), .B2(new_n898_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n899_), .A2(new_n265_), .A3(new_n279_), .A4(new_n283_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1349gat));
  NOR4_X1   g710(.A1(new_n896_), .A2(new_n428_), .A3(new_n349_), .A4(new_n898_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n898_), .A2(new_n349_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n877_), .A2(new_n587_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n404_), .ZN(G1350gat));
  NAND3_X1  g714(.A1(new_n899_), .A2(new_n626_), .A3(new_n438_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n896_), .A2(new_n665_), .A3(new_n898_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n422_), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n897_), .A2(new_n589_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n875_), .A2(new_n876_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n331_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n290_), .A2(KEYINPUT126), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n290_), .A2(KEYINPUT126), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n921_), .B2(new_n923_), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n920_), .A2(new_n884_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G204gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n386_), .B2(new_n926_), .ZN(G1353gat));
  NAND2_X1  g727(.A1(new_n920_), .A2(new_n350_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  XOR2_X1   g729(.A(KEYINPUT63), .B(G211gat), .Z(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(new_n931_), .ZN(G1354gat));
  AOI21_X1  g731(.A(G218gat), .B1(new_n920_), .B2(new_n626_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n919_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n849_), .A2(new_n854_), .A3(G218gat), .A4(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n665_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n933_), .B2(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n849_), .A2(new_n854_), .A3(new_n626_), .A4(new_n934_), .ZN(new_n938_));
  INV_X1    g737(.A(G218gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n940_), .B(new_n941_), .C1(new_n665_), .C2(new_n935_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n937_), .A2(new_n942_), .ZN(G1355gat));
endmodule


