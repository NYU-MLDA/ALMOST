//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G228gat), .A2(G233gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT88), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT29), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR3_X1   g007(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT85), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(KEYINPUT2), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n210_), .B(new_n211_), .C1(new_n222_), .C2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n206_), .B1(new_n219_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT87), .B(G197gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(G204gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n231_), .A2(G204gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(G197gat), .B2(G204gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n234_), .A2(new_n237_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n233_), .A2(new_n239_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n205_), .B1(new_n229_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(new_n240_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n231_), .A2(G204gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n238_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n234_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n204_), .B(KEYINPUT88), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n220_), .B(KEYINPUT85), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n250_), .A2(new_n225_), .A3(new_n226_), .A4(new_n223_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n208_), .A2(new_n209_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(G155gat), .B2(G162gat), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n251_), .A2(new_n253_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n248_), .B(new_n249_), .C1(new_n254_), .C2(new_n206_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n203_), .B1(new_n242_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(KEYINPUT89), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n219_), .A2(new_n228_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT29), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G22gat), .B(G50gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n254_), .A2(new_n206_), .A3(new_n258_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT90), .B1(new_n257_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT90), .ZN(new_n268_));
  OAI221_X1 g067(.A(new_n268_), .B1(new_n264_), .B2(new_n265_), .C1(new_n256_), .C2(KEYINPUT89), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n242_), .A2(new_n255_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(new_n202_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(new_n256_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n267_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT77), .B(G183gat), .Z(new_n279_));
  INV_X1    g078(.A(KEYINPUT25), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT26), .B(G190gat), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT78), .ZN(new_n283_));
  INV_X1    g082(.A(G190gat), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n284_), .A2(KEYINPUT26), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n281_), .B(new_n283_), .C1(KEYINPUT78), .C2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G169gat), .B(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT79), .ZN(new_n290_));
  NOR3_X1   g089(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT79), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n293_), .B(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n298_), .B2(new_n295_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n286_), .A2(new_n290_), .A3(new_n292_), .A4(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G169gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n298_), .A2(new_n295_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n279_), .A2(new_n284_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n303_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G227gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(G15gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT30), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n301_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n301_), .B2(new_n310_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT82), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(KEYINPUT82), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n320_), .A2(KEYINPUT82), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n321_), .A3(new_n318_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT83), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(KEYINPUT83), .A3(new_n326_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n317_), .A2(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n329_), .B(new_n328_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  INV_X1    g133(.A(G43gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT31), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n333_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n277_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G1gat), .B(G29gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT98), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT96), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n324_), .A2(KEYINPUT83), .A3(new_n326_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n260_), .B1(new_n350_), .B2(new_n327_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n254_), .A2(new_n326_), .A3(new_n324_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(KEYINPUT4), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT95), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n351_), .A2(new_n355_), .A3(KEYINPUT4), .A4(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT97), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n351_), .B2(KEYINPUT4), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n330_), .A2(KEYINPUT97), .A3(new_n360_), .A4(new_n260_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n349_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(new_n352_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(new_n348_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n346_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n359_), .A2(new_n361_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n345_), .B(new_n368_), .C1(new_n370_), .C2(new_n349_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n371_), .A3(KEYINPUT100), .ZN(new_n372_));
  XOR2_X1   g171(.A(G8gat), .B(G36gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT32), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT19), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(new_n287_), .B2(new_n384_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n308_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT91), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n282_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n299_), .A2(new_n394_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n388_), .A2(new_n393_), .B1(new_n395_), .B2(new_n303_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n383_), .B1(new_n396_), .B2(new_n241_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n241_), .B1(new_n301_), .B2(new_n310_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n382_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n301_), .A2(new_n241_), .A3(new_n310_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(KEYINPUT20), .C1(new_n396_), .C2(new_n241_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(new_n381_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n379_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT99), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n382_), .A3(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n381_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n378_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT99), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n404_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT100), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n412_), .B(new_n346_), .C1(new_n363_), .C2(new_n366_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n372_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n377_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n303_), .B1(new_n299_), .B2(new_n394_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n387_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n416_), .B1(new_n418_), .B2(new_n392_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT20), .B1(new_n419_), .B2(new_n248_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n420_), .A2(new_n381_), .A3(new_n398_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n383_), .B1(new_n419_), .B2(new_n248_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n382_), .B1(new_n422_), .B2(new_n401_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n415_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n407_), .A2(new_n408_), .A3(new_n377_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n407_), .A2(new_n408_), .A3(KEYINPUT94), .A4(new_n377_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n370_), .A2(new_n349_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n346_), .B1(new_n365_), .B2(new_n348_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n427_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n367_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT33), .B(new_n346_), .C1(new_n363_), .C2(new_n366_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n340_), .B1(new_n414_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n333_), .B(new_n337_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n267_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n273_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n275_), .A2(new_n339_), .A3(new_n276_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n372_), .A2(new_n413_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n427_), .A2(new_n428_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n415_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT27), .A3(new_n425_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n444_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n437_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT6), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  INV_X1    g262(.A(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT9), .A3(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n458_), .A2(new_n462_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n460_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT64), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n471_), .A2(new_n472_), .A3(new_n460_), .A4(KEYINPUT64), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n475_), .A2(new_n458_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n465_), .A2(new_n466_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n470_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  INV_X1    g285(.A(G64gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G57gat), .ZN(new_n488_));
  INV_X1    g287(.A(G57gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G64gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT11), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G71gat), .B(G78gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT66), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(G71gat), .A2(G78gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G71gat), .A2(G78gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n496_), .B(new_n497_), .C1(new_n498_), .C2(KEYINPUT11), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n493_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n493_), .B2(new_n499_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n486_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT11), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n489_), .A2(G64gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n487_), .A2(G57gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n497_), .B1(new_n508_), .B2(new_n496_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n491_), .A2(KEYINPUT66), .A3(new_n492_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n500_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n493_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(KEYINPUT67), .A3(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n485_), .A2(new_n504_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n469_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n470_), .A2(KEYINPUT68), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n478_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n481_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n516_), .B(new_n517_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n514_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n469_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n502_), .A2(new_n503_), .A3(new_n486_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT67), .B1(new_n511_), .B2(new_n512_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n521_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G230gat), .A2(G233gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n514_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G120gat), .B(G148gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n531_), .A2(new_n534_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n541_), .A2(KEYINPUT13), .A3(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(KEYINPUT70), .A3(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  INV_X1    g352(.A(G1gat), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G29gat), .B(G36gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G43gat), .B(G50gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n559_), .B(new_n562_), .Z(new_n563_));
  NAND2_X1  g362(.A1(G229gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n562_), .B(KEYINPUT15), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n559_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n559_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n568_), .B2(new_n562_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n563_), .A2(new_n565_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G113gat), .B(G141gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G169gat), .B(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n570_), .A2(new_n573_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n552_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n453_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT76), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n520_), .B2(new_n566_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n485_), .B2(new_n562_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n562_), .B(new_n469_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT72), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT74), .B(new_n588_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT73), .B(new_n588_), .C1(new_n590_), .C2(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT71), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n584_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n582_), .B(KEYINPUT36), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n593_), .A2(new_n594_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n596_), .A2(new_n598_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n601_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n599_), .A2(KEYINPUT75), .A3(new_n601_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n602_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n607_), .A2(new_n604_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n602_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT37), .ZN(new_n614_));
  OAI22_X1  g413(.A1(new_n611_), .A2(KEYINPUT37), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n559_), .B(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n502_), .A2(new_n503_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  OR4_X1    g424(.A1(new_n616_), .A2(new_n620_), .A3(new_n621_), .A4(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n504_), .A2(new_n513_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n627_), .B1(new_n618_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n618_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n579_), .B1(new_n615_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n612_), .A2(new_n633_), .A3(new_n602_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n607_), .A2(new_n608_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n610_), .A3(new_n603_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n613_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n637_), .B2(new_n633_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n631_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(KEYINPUT76), .A3(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n578_), .A2(new_n632_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n444_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n554_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n631_), .B(new_n611_), .C1(new_n437_), .C2(new_n452_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n577_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n444_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n644_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n648_), .A3(new_n649_), .ZN(G1324gat));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n555_), .A3(new_n450_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n647_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n555_), .B1(new_n652_), .B2(new_n450_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n653_), .A2(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n651_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1325gat));
  NAND3_X1  g459(.A1(new_n641_), .A2(new_n312_), .A3(new_n438_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT102), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n312_), .B1(new_n652_), .B2(new_n438_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n661_), .A2(KEYINPUT102), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n662_), .A2(new_n665_), .A3(new_n666_), .A4(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n647_), .B2(new_n277_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n277_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n641_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n611_), .A2(new_n631_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT105), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n578_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(G29gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(new_n642_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n577_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n639_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n443_), .A2(new_n444_), .A3(new_n451_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n615_), .B1(new_n682_), .B2(new_n436_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT43), .B1(new_n683_), .B2(KEYINPUT103), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n681_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n642_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n688_), .A2(KEYINPUT104), .A3(new_n642_), .A4(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G29gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n679_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT106), .B(new_n679_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1328gat));
  NOR2_X1   g498(.A1(new_n451_), .A2(G36gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n677_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT45), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n677_), .A2(new_n703_), .A3(new_n700_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n702_), .A2(new_n704_), .B1(KEYINPUT107), .B2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n688_), .A2(new_n450_), .A3(new_n689_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G36gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1329gat));
  NOR2_X1   g510(.A1(new_n339_), .A2(new_n335_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n688_), .A2(new_n689_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n688_), .A2(KEYINPUT108), .A3(new_n689_), .A4(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G43gat), .B1(new_n677_), .B2(new_n438_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT109), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n717_), .A2(new_n722_), .A3(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1330gat));
  INV_X1    g523(.A(G50gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n677_), .A2(new_n725_), .A3(new_n672_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n688_), .A2(new_n672_), .A3(new_n689_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT110), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n688_), .A2(new_n729_), .A3(new_n672_), .A4(new_n689_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT111), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n726_), .C1(new_n728_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1331gat));
  INV_X1    g535(.A(new_n552_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n576_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n453_), .A2(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(new_n632_), .A3(new_n640_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n489_), .A3(new_n642_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n646_), .A2(new_n739_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n444_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1332gat));
  OAI21_X1  g544(.A(G64gat), .B1(new_n743_), .B2(new_n451_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT48), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n487_), .A3(new_n450_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1333gat));
  OAI21_X1  g548(.A(G71gat), .B1(new_n743_), .B2(new_n339_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT49), .ZN(new_n751_));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n752_), .A3(new_n438_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n743_), .B2(new_n277_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n741_), .A2(new_n757_), .A3(new_n672_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1335gat));
  OR2_X1    g558(.A1(new_n684_), .A2(new_n685_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n737_), .A2(new_n639_), .A3(new_n738_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n444_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n740_), .A2(new_n676_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n463_), .A3(new_n642_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1336gat));
  NAND2_X1  g565(.A1(new_n450_), .A2(G92gat), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT113), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n760_), .A2(new_n761_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n764_), .A2(new_n450_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n464_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT112), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT112), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT114), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n769_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n762_), .B2(new_n339_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n764_), .A2(new_n459_), .A3(new_n461_), .A4(new_n438_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n764_), .A2(new_n460_), .A3(new_n672_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n761_), .B(new_n672_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g589(.A1(new_n444_), .A2(new_n450_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n441_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n738_), .A2(new_n543_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n483_), .A2(new_n484_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n504_), .A2(new_n513_), .B1(new_n797_), .B2(new_n469_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n514_), .B(new_n523_), .C1(new_n798_), .C2(KEYINPUT12), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n799_), .B2(new_n533_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n533_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n524_), .A2(new_n529_), .A3(KEYINPUT55), .A4(new_n530_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n540_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n530_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n531_), .B1(new_n808_), .B2(new_n796_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n803_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n540_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n795_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n564_), .B1(new_n568_), .B2(new_n562_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n567_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n573_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n574_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n544_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT57), .B(new_n637_), .C1(new_n812_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n637_), .B1(new_n812_), .B2(new_n818_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n795_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n540_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n806_), .B(new_n542_), .C1(new_n809_), .C2(new_n803_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n817_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n637_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n816_), .A2(new_n543_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n831_), .B(KEYINPUT58), .C1(new_n826_), .C2(new_n827_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n615_), .A3(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n821_), .A2(new_n824_), .A3(new_n830_), .A4(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n631_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NAND2_X1  g638(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n631_), .A2(new_n738_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n546_), .A2(new_n547_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n843_), .B1(new_n638_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT37), .B1(new_n636_), .B2(new_n613_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n848_), .A2(new_n845_), .A3(new_n634_), .A4(new_n841_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n839_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n615_), .A2(new_n845_), .B1(new_n842_), .B2(new_n841_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n638_), .A2(new_n846_), .A3(new_n840_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(KEYINPUT117), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n838_), .A2(new_n854_), .A3(KEYINPUT119), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT119), .B1(new_n838_), .B2(new_n854_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n794_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n738_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n838_), .A2(new_n854_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n793_), .A2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n860_), .B1(new_n861_), .B2(new_n866_), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT121), .B(new_n865_), .C1(new_n857_), .C2(KEYINPUT59), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n738_), .A2(G113gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n859_), .B1(new_n869_), .B2(new_n870_), .ZN(G1340gat));
  AOI211_X1 g670(.A(new_n737_), .B(new_n865_), .C1(new_n857_), .C2(KEYINPUT59), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT122), .B(G120gat), .Z(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT123), .B1(new_n873_), .B2(KEYINPUT60), .ZN(new_n874_));
  INV_X1    g673(.A(new_n873_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n552_), .B2(new_n876_), .ZN(new_n877_));
  MUX2_X1   g676(.A(new_n874_), .B(KEYINPUT123), .S(new_n877_), .Z(new_n878_));
  OAI22_X1  g677(.A1(new_n872_), .A2(new_n873_), .B1(new_n857_), .B2(new_n878_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n858_), .B2(new_n639_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n639_), .A2(G127gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n869_), .B2(new_n882_), .ZN(G1342gat));
  AOI21_X1  g682(.A(G134gat), .B1(new_n858_), .B2(new_n611_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n615_), .A2(G134gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n869_), .B2(new_n885_), .ZN(G1343gat));
  OR2_X1    g685(.A1(new_n855_), .A2(new_n856_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n444_), .A2(new_n442_), .A3(new_n450_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n738_), .A3(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n552_), .A3(new_n888_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  OAI211_X1 g691(.A(new_n639_), .B(new_n888_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n893_), .A2(KEYINPUT124), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(KEYINPUT124), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1346gat));
  NAND2_X1  g698(.A1(new_n887_), .A2(new_n888_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G162gat), .B1(new_n900_), .B2(new_n638_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n637_), .A2(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(new_n902_), .ZN(G1347gat));
  NAND3_X1  g702(.A1(new_n444_), .A2(new_n438_), .A3(new_n450_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n672_), .B(new_n904_), .C1(new_n838_), .C2(new_n854_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n738_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906_), .B2(KEYINPUT62), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT62), .B1(new_n906_), .B2(KEYINPUT22), .ZN(new_n908_));
  MUX2_X1   g707(.A(G169gat), .B(new_n907_), .S(new_n908_), .Z(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n905_), .B2(new_n552_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n887_), .A2(new_n277_), .ZN(new_n911_));
  INV_X1    g710(.A(G176gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n737_), .A2(new_n912_), .A3(new_n904_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n911_), .B2(new_n913_), .ZN(G1349gat));
  NOR2_X1   g713(.A1(new_n904_), .A2(new_n631_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n639_), .A2(new_n391_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n916_), .A2(new_n279_), .B1(new_n905_), .B2(new_n918_), .ZN(G1350gat));
  NOR2_X1   g718(.A1(new_n637_), .A2(new_n282_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n905_), .A2(new_n920_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n905_), .A2(new_n615_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n284_), .ZN(G1351gat));
  NAND3_X1  g722(.A1(new_n444_), .A2(new_n672_), .A3(new_n339_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n450_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n925_), .B2(new_n924_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(KEYINPUT126), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT126), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n930_), .B(new_n927_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n576_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(G197gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1352gat));
  AOI21_X1  g733(.A(new_n737_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n935_));
  INV_X1    g734(.A(G204gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1353gat));
  OR3_X1    g736(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n639_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n941_), .B(new_n942_), .ZN(G1354gat));
  NAND2_X1  g742(.A1(new_n929_), .A2(new_n931_), .ZN(new_n944_));
  INV_X1    g743(.A(G218gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(new_n945_), .A3(new_n611_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n638_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n945_), .ZN(G1355gat));
endmodule


