//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n204_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(G92gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n210_), .A2(new_n215_), .A3(new_n218_), .A4(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n213_), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT66), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n212_), .A2(new_n214_), .A3(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(new_n227_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n222_), .B1(new_n232_), .B2(new_n219_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n219_), .A2(new_n222_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n234_), .B1(new_n215_), .B2(new_n231_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n221_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G57gat), .B(G64gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(KEYINPUT11), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n239_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n243_), .B(new_n221_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n248_), .A3(new_n244_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n203_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n202_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G120gat), .B(G148gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G176gat), .B(G204gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT67), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n252_), .A2(new_n259_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263_));
  OAI22_X1  g062(.A1(new_n261_), .A2(new_n262_), .B1(new_n263_), .B2(KEYINPUT13), .ZN(new_n264_));
  INV_X1    g063(.A(new_n262_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n260_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n268_), .A2(KEYINPUT69), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(KEYINPUT69), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G43gat), .B(G50gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G36gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G29gat), .ZN(new_n276_));
  INV_X1    g075(.A(G29gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G36gat), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT70), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT70), .B1(new_n276_), .B2(new_n278_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n274_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n278_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n276_), .A2(new_n278_), .A3(KEYINPUT70), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n285_), .A3(new_n273_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n287_), .B(new_n221_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT71), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G232gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT34), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT35), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT72), .B1(new_n291_), .B2(KEYINPUT35), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n281_), .A2(new_n286_), .A3(KEYINPUT15), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT15), .B1(new_n281_), .B2(new_n286_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(new_n236_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n289_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n292_), .B1(new_n289_), .B2(new_n297_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G190gat), .B(G218gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G134gat), .B(G162gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT36), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n303_), .A2(KEYINPUT36), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n300_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n289_), .A2(new_n297_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n292_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n289_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(KEYINPUT73), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n272_), .B(new_n305_), .C1(new_n308_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT37), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n300_), .A2(new_n304_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(KEYINPUT73), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n300_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n321_), .A2(new_n272_), .A3(KEYINPUT37), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G231gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT76), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n243_), .B(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G1gat), .A2(G8gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G1gat), .A2(G8gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(new_n332_), .B2(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G15gat), .B(G22gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n330_), .A2(KEYINPUT14), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n331_), .A2(new_n333_), .A3(new_n336_), .A4(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n326_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G127gat), .B(G155gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT16), .ZN(new_n343_));
  XOR2_X1   g142(.A(G183gat), .B(G211gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT17), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT17), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n341_), .B1(new_n348_), .B2(new_n345_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n271_), .A2(new_n323_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT77), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(G169gat), .B2(G176gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G183gat), .A2(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n354_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G190gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT25), .B(G183gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n357_), .B(new_n358_), .C1(G183gat), .C2(G190gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G169gat), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n361_), .A2(new_n364_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT30), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  INV_X1    g169(.A(G15gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G71gat), .ZN(new_n373_));
  INV_X1    g172(.A(G99gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n369_), .A2(new_n375_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G127gat), .B(G134gat), .Z(new_n379_));
  XOR2_X1   g178(.A(G113gat), .B(G120gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT31), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n376_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n383_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT80), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G141gat), .ZN(new_n395_));
  INV_X1    g194(.A(G148gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT81), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT2), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT3), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(G141gat), .B2(G148gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT2), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT81), .B(new_n404_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n404_), .A2(new_n410_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT82), .A3(new_n398_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n394_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n393_), .B(KEYINPUT1), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n392_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G141gat), .B(G148gat), .Z(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n381_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n394_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT82), .B1(new_n411_), .B2(new_n398_), .ZN(new_n423_));
  AND4_X1   g222(.A1(KEYINPUT82), .A2(new_n398_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n381_), .A3(new_n417_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT92), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT83), .B1(new_n413_), .B2(new_n418_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n430_), .A3(new_n417_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n431_), .A3(new_n382_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n429_), .A2(new_n431_), .A3(KEYINPUT91), .A4(new_n382_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n428_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G1gat), .B(G29gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G85gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT0), .B(G57gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n440_), .B(new_n441_), .Z(new_n442_));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443_));
  AOI211_X1 g242(.A(new_n443_), .B(new_n428_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n437_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n432_), .B2(KEYINPUT4), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n438_), .B(new_n442_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n442_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(new_n448_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n438_), .B(new_n451_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G8gat), .B(G36gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT18), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G226gat), .A2(G233gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G211gat), .B(G218gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT21), .ZN(new_n464_));
  AND2_X1   g263(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(KEYINPUT86), .A2(G204gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(G197gat), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G197gat), .A2(G204gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT87), .B1(new_n464_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT86), .B(G204gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n468_), .B1(new_n472_), .B2(G197gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT21), .A4(new_n463_), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n465_), .A2(new_n466_), .A3(G197gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT21), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(G197gat), .B2(G204gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n463_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n477_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n471_), .A2(new_n475_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT89), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n363_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n363_), .A2(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n362_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n485_), .A2(new_n361_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT20), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n471_), .A2(new_n475_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n479_), .A2(new_n480_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n488_), .A2(new_n368_), .A3(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n458_), .B(new_n462_), .C1(new_n487_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n489_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n368_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n496_), .A3(new_n461_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n481_), .A2(new_n368_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(KEYINPUT20), .C1(new_n481_), .C2(new_n486_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n458_), .B1(new_n500_), .B2(new_n462_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n457_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n462_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT90), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(new_n456_), .A3(new_n497_), .A4(new_n491_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n436_), .A2(KEYINPUT4), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n432_), .A2(KEYINPUT4), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(new_n445_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n442_), .B1(new_n436_), .B2(new_n445_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n506_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n449_), .A2(new_n452_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n446_), .B1(new_n436_), .B2(KEYINPUT4), .ZN(new_n514_));
  AOI211_X1 g313(.A(new_n445_), .B(new_n428_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n450_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n447_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n461_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n518_), .A2(new_n519_), .B1(new_n500_), .B2(new_n462_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n518_), .A2(new_n519_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT32), .B(new_n456_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n456_), .A2(KEYINPUT32), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n504_), .A2(new_n497_), .A3(new_n491_), .A4(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n429_), .A2(new_n431_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT28), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT84), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT28), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n528_), .A2(new_n533_), .A3(new_n529_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n536_));
  AOI211_X1 g335(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n429_), .C2(new_n431_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT84), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G22gat), .B(G50gat), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n429_), .A2(new_n431_), .A3(KEYINPUT29), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G228gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n481_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n494_), .B1(new_n419_), .B2(new_n529_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n542_), .A2(new_n545_), .B1(new_n546_), .B2(new_n544_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G78gat), .B(G106gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT85), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n540_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n535_), .A2(new_n538_), .A3(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n541_), .A2(new_n549_), .A3(new_n551_), .A4(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n551_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n535_), .A2(new_n538_), .A3(new_n552_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n552_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n513_), .A2(new_n527_), .B1(new_n554_), .B2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n505_), .A2(KEYINPUT27), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n457_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT94), .B(KEYINPUT27), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n560_), .A2(new_n561_), .B1(new_n506_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n564_), .A2(new_n517_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n390_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n554_), .A2(new_n558_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n563_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n517_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n389_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n340_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n287_), .A2(new_n339_), .A3(new_n338_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n281_), .A2(new_n286_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n340_), .A2(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n338_), .A2(new_n339_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(KEYINPUT78), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n575_), .A2(new_n585_), .A3(new_n576_), .A4(new_n577_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n586_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n573_), .A2(new_n574_), .A3(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n569_), .A2(new_n554_), .A3(new_n558_), .A4(new_n563_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n525_), .B1(new_n516_), .B2(new_n447_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n510_), .A2(new_n511_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n506_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n598_), .A2(new_n452_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n597_), .B1(new_n600_), .B2(new_n449_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n567_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n596_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n571_), .B1(new_n603_), .B2(new_n390_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n584_), .A2(new_n586_), .A3(new_n592_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n592_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT95), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n352_), .B1(new_n595_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(G1gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n517_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n321_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n573_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n268_), .A2(new_n594_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n350_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n569_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n611_), .A2(new_n612_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n613_), .A2(new_n621_), .A3(new_n622_), .ZN(G1324gat));
  INV_X1    g422(.A(G8gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n563_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n609_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n616_), .A2(new_n625_), .A3(new_n619_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(new_n628_), .A3(G8gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(G8gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n620_), .B2(new_n390_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT96), .B(KEYINPUT41), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT97), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n636_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n609_), .A2(new_n371_), .A3(new_n389_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(G1326gat));
  OAI21_X1  g439(.A(G22gat), .B1(new_n620_), .B2(new_n567_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT42), .ZN(new_n642_));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n609_), .A2(new_n643_), .A3(new_n602_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n608_), .A2(new_n595_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n614_), .A2(new_n350_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n268_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G29gat), .B1(new_n651_), .B2(new_n517_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n604_), .B2(new_n323_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n317_), .A2(new_n322_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n573_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n617_), .A2(new_n350_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(new_n658_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n660_), .B(new_n661_), .C1(new_n653_), .C2(new_n656_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n569_), .A2(new_n277_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n652_), .B1(new_n663_), .B2(new_n664_), .ZN(G1328gat));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT98), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT99), .Z(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n563_), .A2(G36gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n574_), .B1(new_n573_), .B2(new_n594_), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT95), .B(new_n607_), .C1(new_n566_), .C2(new_n572_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n650_), .B(new_n670_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n646_), .A2(KEYINPUT45), .A3(new_n650_), .A4(new_n670_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n654_), .B1(new_n573_), .B2(new_n655_), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT43), .B(new_n323_), .C1(new_n566_), .C2(new_n572_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n660_), .B1(new_n680_), .B2(new_n661_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n657_), .A2(KEYINPUT44), .A3(new_n658_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n625_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n677_), .B1(new_n683_), .B2(G36gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n666_), .A2(KEYINPUT98), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n669_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n685_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n275_), .B1(new_n663_), .B2(new_n625_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n687_), .B(new_n668_), .C1(new_n688_), .C2(new_n677_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(G1329gat));
  NAND4_X1  g489(.A1(new_n681_), .A2(G43gat), .A3(new_n389_), .A4(new_n682_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n646_), .A2(new_n389_), .A3(new_n650_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n693_));
  INV_X1    g492(.A(G43gat), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g497(.A(G50gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n651_), .A2(new_n699_), .A3(new_n602_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n663_), .A2(new_n701_), .A3(new_n602_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n663_), .B2(new_n602_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  NAND2_X1  g504(.A1(new_n350_), .A2(new_n607_), .ZN(new_n706_));
  OR4_X1    g505(.A1(new_n604_), .A2(new_n321_), .A3(new_n271_), .A4(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n569_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n604_), .A2(new_n594_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n710_), .A2(new_n350_), .A3(new_n323_), .A4(new_n649_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n569_), .B1(new_n713_), .B2(KEYINPUT103), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(KEYINPUT103), .B2(new_n713_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n709_), .B1(new_n715_), .B2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n707_), .B2(new_n563_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT48), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n563_), .A2(G64gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n713_), .B2(new_n719_), .ZN(G1333gat));
  XNOR2_X1  g519(.A(new_n711_), .B(KEYINPUT102), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n390_), .A2(G71gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n271_), .A2(new_n706_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n616_), .A2(new_n389_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G71gat), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT49), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT104), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n723_), .B(new_n731_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n707_), .B2(new_n567_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n567_), .A2(G78gat), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT105), .Z(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n713_), .B2(new_n737_), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n271_), .A2(new_n648_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n710_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT106), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n710_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n517_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(KEYINPUT107), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(KEYINPUT107), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n649_), .A2(new_n607_), .A3(new_n618_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT108), .Z(new_n750_));
  AND2_X1   g549(.A1(new_n517_), .A2(new_n216_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n746_), .A2(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  INV_X1    g551(.A(G92gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n744_), .A2(new_n753_), .A3(new_n625_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n750_), .A2(new_n625_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n753_), .ZN(G1337gat));
  OAI21_X1  g555(.A(new_n389_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n744_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n749_), .A2(new_n389_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G99gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n757_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n374_), .B1(new_n749_), .B2(new_n389_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n763_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1338gat));
  NAND3_X1  g569(.A1(new_n744_), .A2(new_n204_), .A3(new_n602_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n749_), .A2(new_n602_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(G106gat), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT52), .B(new_n204_), .C1(new_n749_), .C2(new_n602_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(KEYINPUT112), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n706_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n317_), .A2(new_n322_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(KEYINPUT112), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n317_), .A2(new_n322_), .A3(new_n781_), .A4(new_n783_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n780_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n250_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n607_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n247_), .A2(new_n249_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n202_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n251_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n257_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n594_), .A2(new_n794_), .A3(KEYINPUT113), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n790_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n247_), .A2(new_n203_), .A3(new_n249_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT114), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n247_), .A2(new_n800_), .A3(new_n203_), .A4(new_n249_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n250_), .A2(KEYINPUT55), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n203_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n797_), .B1(new_n806_), .B2(new_n257_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n792_), .A2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n250_), .A2(KEYINPUT55), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n799_), .A4(new_n801_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n256_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n796_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n261_), .A2(new_n262_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n581_), .A2(new_n582_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n576_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n575_), .A2(new_n579_), .A3(new_n577_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n592_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n591_), .A2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n614_), .B1(new_n812_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n607_), .A2(new_n789_), .A3(new_n788_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT113), .B1(new_n594_), .B2(new_n794_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n256_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n256_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n813_), .A2(new_n818_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n614_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n818_), .A2(new_n789_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n811_), .B1(new_n827_), .B2(KEYINPUT115), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n803_), .A2(new_n805_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n799_), .A2(new_n801_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n257_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(KEYINPUT56), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT58), .B(new_n832_), .C1(new_n833_), .C2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n655_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n836_), .B2(KEYINPUT56), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n827_), .A2(KEYINPUT115), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n811_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT58), .B1(new_n843_), .B2(new_n832_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n822_), .B(new_n831_), .C1(new_n840_), .C2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n787_), .B1(new_n845_), .B2(new_n618_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n568_), .A2(new_n569_), .A3(new_n390_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n778_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n614_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n821_), .B(new_n321_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n832_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n655_), .A3(new_n839_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n350_), .B1(new_n852_), .B2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT59), .B(new_n847_), .C1(new_n857_), .C2(new_n787_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n849_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n849_), .A2(KEYINPUT116), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863_), .B2(new_n607_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n846_), .A2(new_n848_), .ZN(new_n865_));
  INV_X1    g664(.A(G113gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n594_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n268_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n865_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n869_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n271_), .B1(new_n849_), .B2(new_n858_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1341gat));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n849_), .A2(KEYINPUT116), .A3(new_n858_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT116), .B1(new_n849_), .B2(new_n858_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n350_), .A2(G127gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n846_), .A2(new_n618_), .A3(new_n848_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(G127gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n874_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n880_), .ZN(new_n882_));
  OAI211_X1 g681(.A(KEYINPUT117), .B(new_n882_), .C1(new_n863_), .C2(new_n877_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1342gat));
  XOR2_X1   g683(.A(KEYINPUT118), .B(G134gat), .Z(new_n885_));
  NOR3_X1   g684(.A1(new_n863_), .A2(new_n323_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G134gat), .B1(new_n865_), .B2(new_n321_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1343gat));
  INV_X1    g687(.A(new_n846_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n564_), .A2(new_n569_), .A3(new_n389_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT119), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n607_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n395_), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n271_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT120), .B(G148gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n892_), .A2(new_n618_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n892_), .B2(new_n323_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n614_), .A2(G162gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n892_), .B2(new_n902_), .ZN(G1347gat));
  XNOR2_X1  g702(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(KEYINPUT123), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n567_), .A2(new_n625_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n570_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n846_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n594_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT121), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n913_), .A3(new_n594_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(G169gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n905_), .B2(KEYINPUT123), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n906_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n906_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n917_), .ZN(new_n920_));
  AOI211_X1 g719(.A(new_n919_), .B(new_n920_), .C1(new_n912_), .C2(new_n914_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT22), .B(G169gat), .Z(new_n922_));
  OAI22_X1  g721(.A1(new_n918_), .A2(new_n921_), .B1(new_n911_), .B2(new_n922_), .ZN(G1348gat));
  INV_X1    g722(.A(new_n910_), .ZN(new_n924_));
  OR3_X1    g723(.A1(new_n924_), .A2(G176gat), .A3(new_n268_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G176gat), .B1(new_n924_), .B2(new_n271_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1349gat));
  AOI21_X1  g726(.A(G183gat), .B1(new_n910_), .B2(new_n350_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n924_), .A2(new_n618_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n483_), .A2(new_n484_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT124), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n910_), .A2(new_n362_), .A3(new_n321_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n910_), .A2(new_n655_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n934_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n935_));
  AOI21_X1  g734(.A(KEYINPUT125), .B1(new_n934_), .B2(G190gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n933_), .B1(new_n935_), .B2(new_n936_), .ZN(G1351gat));
  NAND4_X1  g736(.A1(new_n602_), .A2(new_n569_), .A3(new_n625_), .A4(new_n390_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n846_), .A2(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT126), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n594_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g741(.A(new_n271_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(G204gat), .ZN(new_n945_));
  AND4_X1   g744(.A1(new_n472_), .A2(new_n940_), .A3(new_n943_), .A4(new_n945_), .ZN(new_n946_));
  AOI22_X1  g745(.A1(new_n940_), .A2(new_n943_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1353gat));
  OR2_X1    g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  NAND2_X1  g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  AND4_X1   g749(.A1(new_n350_), .A2(new_n940_), .A3(new_n949_), .A4(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n940_), .B2(new_n350_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1354gat));
  INV_X1    g752(.A(G218gat), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n940_), .A2(new_n954_), .A3(new_n321_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n940_), .A2(new_n655_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n954_), .ZN(G1355gat));
endmodule


