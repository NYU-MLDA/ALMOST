//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G197gat), .ZN(new_n211_));
  INV_X1    g010(.A(G197gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G204gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n209_), .A2(KEYINPUT90), .A3(new_n214_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n210_), .A2(G197gat), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n214_), .B(KEYINPUT21), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n207_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT21), .B1(new_n220_), .B2(new_n219_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n211_), .A2(new_n213_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n217_), .A2(new_n218_), .B1(new_n221_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT95), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT94), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(KEYINPUT22), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT94), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(G176gat), .B1(new_n232_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT93), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n227_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G176gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n236_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n235_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n239_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT95), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT23), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(G183gat), .A3(G190gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT82), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G183gat), .ZN(new_n251_));
  INV_X1    g050(.A(G190gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT23), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n247_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n240_), .A2(new_n246_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G190gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT92), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n228_), .A2(new_n241_), .A3(KEYINPUT81), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT81), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(G169gat), .B2(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n238_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n253_), .A2(new_n248_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(new_n228_), .A3(new_n241_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n261_), .A2(new_n266_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n226_), .B1(new_n257_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n262_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n260_), .A2(new_n258_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n266_), .A2(new_n255_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n234_), .A2(KEYINPUT83), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT83), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n228_), .A3(KEYINPUT22), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n275_), .A2(new_n277_), .A3(new_n241_), .A4(new_n233_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n253_), .A2(new_n248_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n238_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n274_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n223_), .A2(new_n224_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n221_), .A2(new_n284_), .A3(new_n207_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT90), .B1(new_n209_), .B2(new_n214_), .ZN(new_n286_));
  NOR4_X1   g085(.A1(new_n224_), .A2(new_n207_), .A3(new_n216_), .A4(new_n208_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n206_), .B1(new_n271_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n257_), .A2(new_n226_), .A3(new_n270_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT20), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(new_n283_), .B2(new_n288_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n205_), .A3(new_n299_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n290_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n296_), .B1(new_n290_), .B2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n202_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n271_), .A2(new_n206_), .A3(new_n289_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n205_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n295_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n290_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT99), .A4(KEYINPUT27), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(KEYINPUT27), .A3(new_n307_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT99), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G228gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT88), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT86), .B1(new_n318_), .B2(KEYINPUT1), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(G155gat), .A4(G162gat), .ZN(new_n322_));
  INV_X1    g121(.A(G155gat), .ZN(new_n323_));
  INV_X1    g122(.A(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n319_), .A2(new_n322_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G141gat), .B(G148gat), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330_));
  INV_X1    g129(.A(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G148gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n325_), .A2(new_n318_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n288_), .B(new_n316_), .C1(new_n317_), .C2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n329_), .A2(new_n340_), .A3(KEYINPUT87), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n226_), .B1(new_n347_), .B2(KEYINPUT29), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n348_), .B2(new_n316_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(KEYINPUT29), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI221_X1 g150(.A(new_n343_), .B1(KEYINPUT29), .B2(new_n347_), .C1(new_n348_), .C2(new_n316_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G22gat), .B(G50gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT28), .ZN(new_n354_));
  XOR2_X1   g153(.A(G78gat), .B(G106gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n351_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  INV_X1    g161(.A(G113gat), .ZN(new_n363_));
  INV_X1    g162(.A(G120gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G113gat), .A2(G120gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT85), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n369_), .A3(new_n366_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n342_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n372_), .A2(new_n373_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n329_), .A2(new_n340_), .A3(KEYINPUT87), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT87), .B1(new_n329_), .B2(new_n340_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n362_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT4), .B1(new_n347_), .B2(new_n376_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n361_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n379_), .A3(new_n360_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G227gat), .ZN(new_n393_));
  INV_X1    g192(.A(G233gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n376_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n376_), .A2(new_n395_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT30), .B(G15gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n398_), .B(KEYINPUT31), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n396_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G71gat), .B(G99gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G43gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n283_), .B(new_n404_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n401_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n359_), .A2(new_n392_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT101), .B1(new_n313_), .B2(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n312_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT101), .ZN(new_n412_));
  INV_X1    g211(.A(new_n358_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n351_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(new_n412_), .A3(new_n392_), .A4(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n410_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT100), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT32), .B(new_n296_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n296_), .A2(KEYINPUT32), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n290_), .A2(new_n300_), .A3(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n420_), .B(new_n422_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n375_), .A2(new_n379_), .A3(new_n361_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n387_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT97), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT97), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n427_), .A3(new_n387_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n360_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n426_), .A2(new_n429_), .A3(KEYINPUT98), .A4(new_n428_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n382_), .A2(KEYINPUT33), .A3(new_n383_), .A4(new_n388_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n301_), .A2(new_n302_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n389_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n423_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n391_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n389_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n359_), .A2(new_n442_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n359_), .A2(new_n440_), .B1(new_n411_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n419_), .B1(new_n444_), .B2(new_n408_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n359_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n408_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(KEYINPUT100), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n418_), .B1(new_n445_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n452_));
  AND2_X1   g251(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n460_), .A2(KEYINPUT10), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(KEYINPUT10), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT10), .B(G99gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT64), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT65), .B(G106gat), .Z(new_n467_));
  AOI21_X1  g266(.A(new_n458_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT67), .ZN(new_n469_));
  OR2_X1    g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G85gat), .A2(G92gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n470_), .B1(new_n473_), .B2(KEYINPUT9), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT9), .ZN(new_n475_));
  AND2_X1   g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n478_), .B2(new_n471_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n469_), .B1(new_n474_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(KEYINPUT9), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT67), .A4(new_n470_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n468_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n460_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n478_), .B1(new_n489_), .B2(new_n458_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT8), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n484_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT68), .B(G71gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(G78gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G57gat), .B(G64gat), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(G78gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G78gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n493_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n495_), .B(KEYINPUT11), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n498_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n453_), .B1(new_n492_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n484_), .A2(new_n491_), .A3(new_n502_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n502_), .B1(new_n484_), .B2(new_n491_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n453_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n510_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n505_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n511_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n210_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT5), .B(G176gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n452_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n513_), .A2(new_n516_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n520_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n521_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532_));
  INV_X1    g331(.A(G50gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(G43gat), .ZN(new_n534_));
  INV_X1    g333(.A(G43gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G50gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n539_));
  INV_X1    g338(.A(G36gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G29gat), .ZN(new_n541_));
  INV_X1    g340(.A(G29gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G36gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n538_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n541_), .A2(new_n543_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n535_), .A2(G50gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n533_), .A2(G43gat), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT71), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n532_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n544_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n550_), .A3(new_n546_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT15), .ZN(new_n555_));
  XOR2_X1   g354(.A(G15gat), .B(G22gat), .Z(new_n556_));
  OR2_X1    g355(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(G8gat), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n556_), .B1(KEYINPUT14), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G1gat), .B(G8gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT75), .ZN(new_n562_));
  OR2_X1    g361(.A1(G1gat), .A2(G8gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G1gat), .A2(G8gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n566_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n559_), .A2(KEYINPUT14), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n569_), .B2(new_n556_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n552_), .A2(new_n555_), .A3(new_n567_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT78), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G229gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n560_), .B(new_n568_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT78), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n555_), .A4(new_n552_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n545_), .A2(new_n551_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n567_), .A2(new_n570_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n572_), .A2(new_n573_), .A3(new_n576_), .A4(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n573_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n580_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n578_), .A2(new_n579_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT79), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n581_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT80), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  NAND3_X1  g392(.A1(new_n587_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n589_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n588_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n531_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n451_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n552_), .A2(new_n555_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n492_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT34), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT35), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n484_), .A2(new_n491_), .A3(new_n578_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT35), .A3(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(KEYINPUT35), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n605_), .A2(new_n612_), .A3(new_n608_), .A4(new_n609_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(KEYINPUT72), .A3(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n611_), .A2(KEYINPUT72), .A3(new_n619_), .A4(new_n613_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n611_), .A2(new_n613_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n617_), .A2(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n622_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n621_), .A2(new_n625_), .A3(new_n622_), .A4(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n323_), .A2(G127gat), .ZN(new_n633_));
  INV_X1    g432(.A(G127gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G155gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(G211gat), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n635_), .A3(G211gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT16), .B(G183gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n633_), .A2(new_n635_), .A3(G211gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n636_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n640_), .A2(new_n643_), .A3(KEYINPUT17), .ZN(new_n644_));
  INV_X1    g443(.A(G231gat), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n394_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n644_), .A2(KEYINPUT76), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n644_), .B2(KEYINPUT76), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n502_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(KEYINPUT76), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n646_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(KEYINPUT76), .A3(new_n647_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n503_), .A3(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n650_), .A2(new_n654_), .A3(new_n574_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n640_), .A2(new_n643_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT17), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n574_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT77), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT77), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n658_), .A4(new_n655_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n632_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n603_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n392_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT38), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n659_), .A2(new_n660_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n601_), .A2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n626_), .B(KEYINPUT102), .Z(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT103), .B1(new_n451_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n410_), .A2(new_n417_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT100), .B1(new_n448_), .B2(new_n449_), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n419_), .B(new_n408_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n676_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n675_), .B1(new_n678_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G1gat), .B1(new_n686_), .B2(new_n392_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n672_), .A2(new_n687_), .ZN(G1324gat));
  INV_X1    g487(.A(G8gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n669_), .A2(new_n689_), .A3(new_n313_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n685_), .B2(new_n313_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT39), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n691_), .A2(new_n692_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g495(.A(G15gat), .B1(new_n686_), .B2(new_n449_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT41), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(KEYINPUT41), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n668_), .A2(G15gat), .A3(new_n449_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(G1326gat));
  INV_X1    g500(.A(G22gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n359_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n685_), .B2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT42), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n669_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n682_), .A2(new_n632_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n632_), .B2(KEYINPUT104), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n665_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n682_), .A2(new_n632_), .A3(new_n710_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n712_), .A2(KEYINPUT44), .A3(new_n601_), .A4(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n451_), .B2(new_n631_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n715_), .A2(new_n713_), .A3(new_n601_), .A4(new_n666_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n714_), .A2(new_n718_), .A3(new_n442_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n676_), .A2(new_n665_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n603_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n442_), .A2(new_n542_), .ZN(new_n722_));
  OAI22_X1  g521(.A1(new_n719_), .A2(new_n542_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n714_), .A2(new_n718_), .A3(new_n313_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n714_), .A2(new_n718_), .A3(KEYINPUT105), .A4(new_n313_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(G36gat), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n729_));
  NOR2_X1   g528(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n411_), .A2(G36gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n721_), .A2(KEYINPUT45), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT45), .B1(new_n721_), .B2(new_n732_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n728_), .A2(new_n729_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n729_), .B1(new_n728_), .B2(new_n735_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1329gat));
  NOR2_X1   g537(.A1(new_n449_), .A2(new_n535_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n714_), .A2(new_n718_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT107), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n714_), .A2(new_n718_), .A3(new_n742_), .A4(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n535_), .B1(new_n721_), .B2(new_n449_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT47), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1330gat));
  NAND3_X1  g549(.A1(new_n714_), .A2(new_n718_), .A3(new_n703_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G50gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n703_), .A2(new_n533_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT109), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n753_), .A2(new_n754_), .B1(new_n721_), .B2(new_n756_), .ZN(G1331gat));
  NOR2_X1   g556(.A1(new_n530_), .A2(new_n599_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n682_), .A2(new_n667_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n442_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n758_), .ZN(new_n761_));
  AOI211_X1 g560(.A(new_n666_), .B(new_n761_), .C1(new_n678_), .C2(new_n684_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n442_), .A2(G57gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n760_), .B1(new_n762_), .B2(new_n763_), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n411_), .A2(G64gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT110), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(G64gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n762_), .B2(new_n313_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n769_), .A2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(G1333gat));
  INV_X1    g572(.A(G71gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n762_), .B2(new_n408_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n776_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n408_), .A2(new_n774_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT112), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n759_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n777_), .A2(new_n778_), .A3(new_n781_), .ZN(G1334gat));
  NAND3_X1  g581(.A1(new_n759_), .A2(new_n499_), .A3(new_n703_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n499_), .B1(new_n762_), .B2(new_n703_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1335gat));
  AND3_X1   g587(.A1(new_n682_), .A2(new_n720_), .A3(new_n758_), .ZN(new_n789_));
  AOI21_X1  g588(.A(G85gat), .B1(new_n789_), .B2(new_n442_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n715_), .A2(new_n713_), .A3(new_n666_), .A4(new_n758_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n442_), .A2(G85gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(G1336gat));
  AOI21_X1  g593(.A(G92gat), .B1(new_n789_), .B2(new_n313_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n313_), .A2(G92gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n792_), .B2(new_n796_), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n791_), .B2(new_n449_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n789_), .A2(new_n466_), .A3(new_n408_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g600(.A1(new_n789_), .A2(new_n467_), .A3(new_n703_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n712_), .A2(new_n703_), .A3(new_n713_), .A4(new_n758_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n486_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n715_), .A2(new_n713_), .A3(new_n666_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT113), .A3(new_n703_), .A4(new_n758_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n791_), .B2(new_n359_), .ZN(new_n810_));
  AND4_X1   g609(.A1(new_n803_), .A2(new_n808_), .A3(G106gat), .A4(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n802_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n802_), .B(new_n813_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n313_), .A2(new_n392_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n416_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n505_), .B(new_n507_), .C1(new_n511_), .C2(new_n453_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n511_), .A2(new_n453_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n514_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n514_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(KEYINPUT55), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NOR4_X1   g624(.A1(new_n820_), .A2(new_n821_), .A3(new_n825_), .A4(new_n514_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n526_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n510_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n513_), .B1(new_n830_), .B2(new_n825_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n826_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n526_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n572_), .A2(new_n582_), .A3(new_n576_), .A4(new_n580_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n573_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n595_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n594_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n594_), .A2(KEYINPUT119), .A3(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n522_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n835_), .A2(KEYINPUT58), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT58), .B1(new_n835_), .B2(new_n843_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n631_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n596_), .A2(new_n597_), .A3(new_n595_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n593_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n521_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT118), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n599_), .A2(new_n851_), .A3(new_n521_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n526_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n828_), .B(new_n520_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n850_), .B(new_n852_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n527_), .A2(new_n521_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n594_), .A2(KEYINPUT119), .A3(new_n838_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT119), .B1(new_n594_), .B2(new_n838_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT120), .B(new_n856_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n855_), .A2(new_n859_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n676_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(new_n676_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n846_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n673_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT115), .B1(new_n666_), .B2(new_n599_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n665_), .A2(new_n870_), .A3(new_n598_), .A4(new_n594_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n631_), .A2(new_n530_), .A3(new_n869_), .A4(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT117), .B1(new_n872_), .B2(KEYINPUT116), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n869_), .A2(new_n530_), .A3(new_n871_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .A4(new_n631_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT54), .B1(new_n872_), .B2(KEYINPUT116), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n873_), .A2(new_n879_), .A3(new_n877_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n819_), .B1(new_n868_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G113gat), .B1(new_n884_), .B2(new_n599_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n844_), .A2(new_n845_), .A3(new_n631_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n863_), .A2(new_n676_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT57), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n863_), .A2(new_n864_), .A3(new_n676_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n883_), .B1(new_n893_), .B2(new_n674_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n819_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n888_), .A2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n883_), .B1(new_n893_), .B2(new_n665_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n887_), .A3(new_n895_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n600_), .A2(new_n363_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n885_), .B1(new_n901_), .B2(new_n902_), .ZN(G1340gat));
  AOI21_X1  g702(.A(KEYINPUT121), .B1(new_n896_), .B2(KEYINPUT59), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n886_), .B(new_n887_), .C1(new_n894_), .C2(new_n895_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n531_), .B(new_n900_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n898_), .A2(KEYINPUT122), .A3(new_n531_), .A4(new_n900_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(G120gat), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n364_), .B1(new_n530_), .B2(KEYINPUT60), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n884_), .B(new_n911_), .C1(KEYINPUT60), .C2(new_n364_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1341gat));
  AOI21_X1  g712(.A(G127gat), .B1(new_n884_), .B2(new_n665_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT123), .B(G127gat), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n673_), .A2(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n901_), .B2(new_n916_), .ZN(G1342gat));
  AOI21_X1  g716(.A(G134gat), .B1(new_n884_), .B2(new_n677_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n632_), .A2(G134gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n901_), .B2(new_n919_), .ZN(G1343gat));
  AOI21_X1  g719(.A(new_n408_), .B1(new_n868_), .B2(new_n883_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n313_), .A2(new_n392_), .A3(new_n359_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n600_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n331_), .ZN(G1344gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n530_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(KEYINPUT124), .B(G148gat), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1345gat));
  NOR2_X1   g727(.A1(new_n923_), .A2(new_n666_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT61), .B(G155gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1346gat));
  NOR3_X1   g730(.A1(new_n923_), .A2(new_n324_), .A3(new_n631_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n923_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n677_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n324_), .B2(new_n934_), .ZN(G1347gat));
  NAND3_X1  g734(.A1(new_n313_), .A2(new_n392_), .A3(new_n408_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n703_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n899_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n938_), .B(new_n599_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n228_), .B1(new_n938_), .B2(new_n599_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n940_), .A2(new_n941_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n939_), .B1(new_n944_), .B2(new_n945_), .ZN(G1348gat));
  AOI21_X1  g745(.A(G176gat), .B1(new_n938_), .B2(new_n531_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n703_), .B1(new_n868_), .B2(new_n883_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n936_), .A2(new_n241_), .A3(new_n530_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n947_), .B1(new_n948_), .B2(new_n949_), .ZN(G1349gat));
  NOR2_X1   g749(.A1(new_n936_), .A2(new_n666_), .ZN(new_n951_));
  AOI21_X1  g750(.A(G183gat), .B1(new_n948_), .B2(new_n951_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n673_), .A2(new_n260_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n938_), .B2(new_n953_), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n938_), .A2(new_n677_), .A3(new_n259_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n938_), .A2(new_n632_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n252_), .ZN(G1351gat));
  NOR3_X1   g756(.A1(new_n411_), .A2(new_n442_), .A3(new_n359_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n921_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n600_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(new_n212_), .ZN(G1352gat));
  NOR2_X1   g760(.A1(new_n959_), .A2(new_n530_), .ZN(new_n962_));
  XOR2_X1   g761(.A(KEYINPUT126), .B(G204gat), .Z(new_n963_));
  XNOR2_X1  g762(.A(new_n962_), .B(new_n963_), .ZN(G1353gat));
  NAND2_X1  g763(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n674_), .A2(new_n965_), .ZN(new_n966_));
  OR3_X1    g765(.A1(new_n959_), .A2(KEYINPUT127), .A3(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(KEYINPUT127), .B1(new_n959_), .B2(new_n966_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n969_), .B(new_n970_), .ZN(G1354gat));
  AND2_X1   g770(.A1(new_n921_), .A2(new_n958_), .ZN(new_n972_));
  AND3_X1   g771(.A1(new_n972_), .A2(G218gat), .A3(new_n632_), .ZN(new_n973_));
  AOI21_X1  g772(.A(G218gat), .B1(new_n972_), .B2(new_n677_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n973_), .A2(new_n974_), .ZN(G1355gat));
endmodule


