//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n206_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G229gat), .A2(G233gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n219_));
  MUX2_X1   g018(.A(new_n206_), .B(new_n219_), .S(new_n213_), .Z(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n220_), .B2(new_n217_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G113gat), .B(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G197gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n221_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(KEYINPUT99), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT24), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(KEYINPUT79), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n244_), .A2(new_n246_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n238_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n232_), .B(new_n233_), .C1(G183gat), .C2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT80), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT22), .B1(new_n253_), .B2(new_n223_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n235_), .A3(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n252_), .A2(new_n257_), .A3(new_n239_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G120gat), .ZN(new_n262_));
  INV_X1    g061(.A(G127gat), .ZN(new_n263_));
  INV_X1    g062(.A(G134gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G113gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G127gat), .A2(G134gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n262_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G120gat), .A3(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n261_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT31), .B(G43gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n275_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT81), .B(G15gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n279_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G22gat), .B(G50gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n289_));
  INV_X1    g088(.A(G141gat), .ZN(new_n290_));
  INV_X1    g089(.A(G148gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n292_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n303_), .A3(new_n300_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n305_), .A2(new_n293_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n290_), .A2(new_n291_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n302_), .A2(KEYINPUT82), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT82), .B1(new_n302_), .B2(new_n308_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G197gat), .B(G204gat), .Z(new_n316_));
  OR2_X1    g115(.A1(G211gat), .A2(G218gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT21), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G211gat), .A2(G218gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(G211gat), .A2(G218gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G211gat), .A2(G218gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT21), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n316_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n325_), .B(KEYINPUT21), .C1(new_n322_), .C2(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT83), .B(KEYINPUT29), .C1(new_n309_), .C2(new_n310_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n302_), .A2(new_n308_), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n333_), .A2(KEYINPUT84), .A3(new_n312_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT84), .B1(new_n333_), .B2(new_n312_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n327_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(G228gat), .A3(G233gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n313_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n337_), .B(new_n313_), .C1(new_n328_), .C2(new_n331_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT28), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n337_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n312_), .A3(new_n311_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n344_), .B2(new_n339_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n288_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT28), .B1(new_n338_), .B2(new_n340_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n342_), .A3(new_n339_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n287_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT18), .B(G64gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G92gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G169gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n235_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n239_), .A3(new_n252_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n359_));
  NAND2_X1  g158(.A1(KEYINPUT85), .A2(KEYINPUT24), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n236_), .A3(new_n239_), .A4(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n242_), .A2(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n363_));
  AND2_X1   g162(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n362_), .B(new_n363_), .C1(new_n364_), .C2(new_n247_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n361_), .A2(new_n365_), .A3(KEYINPUT86), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT86), .B1(new_n361_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n236_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n232_), .A2(new_n233_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n358_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n324_), .A2(new_n326_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT87), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n259_), .B2(new_n373_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n361_), .A2(new_n365_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n361_), .A2(new_n365_), .A3(KEYINPUT86), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n357_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT87), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n327_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(new_n376_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n381_), .A2(new_n357_), .A3(new_n373_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n327_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n388_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT20), .A4(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT88), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n354_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n354_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n383_), .B1(new_n382_), .B2(new_n327_), .ZN(new_n400_));
  AOI211_X1 g199(.A(KEYINPUT87), .B(new_n373_), .C1(new_n381_), .C2(new_n357_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n392_), .B1(new_n402_), .B2(new_n376_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n398_), .B(new_n399_), .C1(new_n403_), .C2(new_n394_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n396_), .A2(new_n397_), .A3(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT89), .B(new_n354_), .C1(new_n389_), .C2(new_n395_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT98), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT20), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n388_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n399_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n396_), .A2(KEYINPUT27), .A3(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n408_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n409_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n284_), .B(new_n350_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n274_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n333_), .A2(new_n273_), .A3(new_n271_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT93), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(KEYINPUT4), .A3(new_n420_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n425_), .B(new_n274_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n423_), .A2(KEYINPUT90), .A3(new_n424_), .A4(new_n426_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n422_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G85gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G1gat), .B(G29gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT92), .B(G57gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n422_), .A2(new_n429_), .A3(new_n430_), .A4(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT96), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n229_), .B1(new_n417_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n408_), .A2(new_n414_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT98), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n408_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n283_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n442_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(KEYINPUT99), .A3(new_n448_), .A4(new_n350_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT94), .Z(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n412_), .A2(KEYINPUT32), .A3(new_n354_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n441_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n429_), .A2(new_n430_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n456_), .A2(KEYINPUT33), .A3(new_n422_), .A4(new_n437_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n440_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n406_), .B2(new_n405_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n418_), .A2(new_n424_), .A3(new_n420_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n423_), .A2(new_n419_), .A3(new_n426_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n438_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n455_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n346_), .A2(new_n349_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT95), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(new_n448_), .A3(new_n408_), .A4(new_n414_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n405_), .A2(new_n406_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n469_), .A2(new_n464_), .A3(new_n459_), .A4(new_n457_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n455_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n350_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n283_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n450_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT6), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  OR3_X1    g279(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(G85gat), .A2(G92gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT8), .B1(new_n485_), .B2(KEYINPUT68), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n482_), .B(new_n485_), .C1(KEYINPUT68), .C2(KEYINPUT8), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n483_), .A2(KEYINPUT9), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT67), .B(G92gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT66), .B(G85gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n494_));
  AOI211_X1 g293(.A(new_n484_), .B(new_n490_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT10), .B(G99gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(KEYINPUT64), .B(G106gat), .Z(new_n497_));
  OAI21_X1  g296(.A(new_n479_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n488_), .B(new_n489_), .C1(new_n495_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n219_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n206_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT34), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n500_), .B(new_n502_), .C1(KEYINPUT35), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT35), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT74), .B(G134gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G162gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(G190gat), .B(G218gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT36), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT37), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n213_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G57gat), .B(G64gat), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n523_));
  XOR2_X1   g322(.A(G71gat), .B(G78gat), .Z(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n523_), .A2(new_n524_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n520_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT75), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT16), .B(G183gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G211gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(G127gat), .B(G155gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n533_), .B(KEYINPUT17), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT76), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n529_), .A2(new_n535_), .B1(new_n528_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT77), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n518_), .A2(new_n539_), .ZN(new_n540_));
  AOI211_X1 g339(.A(KEYINPUT69), .B(KEYINPUT12), .C1(new_n499_), .C2(new_n527_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT12), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n488_), .A2(new_n489_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n490_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n484_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n498_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n527_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n542_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n541_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n499_), .A2(new_n527_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n547_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G120gat), .B(G148gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT71), .Z(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n554_), .A2(new_n557_), .A3(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n566_), .B(new_n567_), .C1(KEYINPUT72), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT73), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AND4_X1   g374(.A1(new_n228_), .A2(new_n477_), .A3(new_n540_), .A4(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n208_), .A3(new_n442_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT100), .Z(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT38), .ZN(new_n579_));
  INV_X1    g378(.A(new_n517_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n539_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n228_), .A3(new_n573_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n580_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  AOI211_X1 g384(.A(new_n584_), .B(new_n585_), .C1(new_n450_), .C2(new_n476_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n208_), .B1(new_n586_), .B2(new_n442_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT102), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(KEYINPUT38), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n579_), .A2(new_n588_), .A3(new_n589_), .ZN(G1324gat));
  NAND2_X1  g389(.A1(new_n445_), .A2(new_n446_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n576_), .A2(new_n209_), .A3(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT103), .Z(new_n594_));
  AOI21_X1  g393(.A(new_n209_), .B1(new_n586_), .B2(new_n592_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT39), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g397(.A(G15gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n586_), .B2(new_n284_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT104), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT41), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n576_), .A2(new_n599_), .A3(new_n284_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1326gat));
  INV_X1    g403(.A(G22gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n586_), .B2(new_n466_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT42), .Z(new_n607_));
  NAND3_X1  g406(.A1(new_n576_), .A2(new_n605_), .A3(new_n466_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  AND3_X1   g408(.A1(new_n573_), .A2(new_n539_), .A3(new_n228_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n477_), .A2(new_n517_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT105), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(G29gat), .B1(new_n613_), .B2(new_n442_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n477_), .B2(new_n518_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n518_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT43), .B(new_n617_), .C1(new_n450_), .C2(new_n476_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n610_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT44), .B(new_n610_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n614_), .B1(new_n626_), .B2(new_n442_), .ZN(G1328gat));
  INV_X1    g426(.A(KEYINPUT46), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n622_), .A2(new_n624_), .A3(new_n591_), .ZN(new_n629_));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n613_), .A2(new_n630_), .A3(new_n592_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT45), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n632_), .B(KEYINPUT45), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n636_), .B(KEYINPUT46), .C1(new_n630_), .C2(new_n629_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1329gat));
  NAND2_X1  g437(.A1(new_n613_), .A2(new_n284_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n203_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n621_), .A2(G43gat), .A3(new_n284_), .A4(new_n623_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT47), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT47), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n647_), .B(new_n640_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1330gat));
  AOI21_X1  g448(.A(G50gat), .B1(new_n613_), .B2(new_n466_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n350_), .A2(new_n205_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n625_), .B2(new_n651_), .ZN(G1331gat));
  AOI21_X1  g451(.A(new_n228_), .B1(new_n450_), .B2(new_n476_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n574_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n517_), .A3(new_n539_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(G57gat), .A3(new_n442_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT108), .Z(new_n657_));
  INV_X1    g456(.A(new_n540_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n658_), .A2(KEYINPUT107), .A3(new_n573_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT107), .B1(new_n658_), .B2(new_n573_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n653_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G57gat), .B1(new_n661_), .B2(new_n442_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n657_), .A2(new_n662_), .ZN(G1332gat));
  NAND2_X1  g462(.A1(new_n655_), .A2(new_n592_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G64gat), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT109), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(KEYINPUT109), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT48), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n591_), .A2(G64gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT110), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n661_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n672_), .A3(new_n673_), .ZN(G1333gat));
  INV_X1    g473(.A(G71gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n655_), .B2(new_n284_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT49), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n675_), .A3(new_n284_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1334gat));
  INV_X1    g478(.A(G78gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n661_), .A2(new_n680_), .A3(new_n466_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n655_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G78gat), .B1(new_n682_), .B2(new_n350_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT50), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT50), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT111), .B(new_n681_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1335gat));
  NAND4_X1  g489(.A1(new_n653_), .A2(new_n517_), .A3(new_n539_), .A4(new_n574_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n442_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n477_), .A2(new_n518_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT43), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n477_), .A2(new_n615_), .A3(new_n518_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT112), .B1(new_n616_), .B2(new_n618_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n581_), .A2(new_n573_), .A3(new_n228_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n701_), .A2(KEYINPUT113), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(KEYINPUT113), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n448_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n693_), .B1(new_n704_), .B2(new_n492_), .ZN(G1336gat));
  AOI21_X1  g504(.A(G92gat), .B1(new_n692_), .B2(new_n592_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n491_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n708_), .B2(new_n592_), .ZN(G1337gat));
  OR2_X1    g508(.A1(new_n283_), .A2(new_n496_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n691_), .A2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT115), .Z(new_n712_));
  NAND4_X1  g511(.A1(new_n698_), .A2(new_n699_), .A3(new_n284_), .A4(new_n700_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G99gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G99gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT51), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n712_), .B(new_n719_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1338gat));
  OR3_X1    g520(.A1(new_n691_), .A2(new_n497_), .A3(new_n350_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n466_), .B(new_n700_), .C1(new_n616_), .C2(new_n618_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G106gat), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT52), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT52), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g527(.A1(new_n417_), .A2(new_n448_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n215_), .A2(new_n217_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n220_), .B2(new_n217_), .ZN(new_n732_));
  MUX2_X1   g531(.A(new_n732_), .B(new_n221_), .S(new_n225_), .Z(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n568_), .ZN(new_n734_));
  NOR4_X1   g533(.A1(new_n541_), .A2(new_n549_), .A3(new_n556_), .A4(new_n552_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n547_), .A2(new_n548_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT12), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n547_), .A2(new_n548_), .A3(new_n542_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n553_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n556_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n735_), .B1(KEYINPUT55), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n739_), .A2(new_n742_), .A3(new_n556_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n565_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT56), .B(new_n565_), .C1(new_n741_), .C2(new_n743_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(KEYINPUT116), .A3(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n228_), .B(new_n567_), .C1(new_n747_), .C2(KEYINPUT116), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n734_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(KEYINPUT57), .A3(new_n580_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT119), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n221_), .B(new_n227_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n551_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n554_), .B1(new_n754_), .B2(new_n742_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n743_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n745_), .B(new_n564_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n746_), .A2(KEYINPUT116), .A3(new_n747_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n567_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n517_), .B1(new_n761_), .B2(new_n734_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(KEYINPUT57), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n746_), .A2(new_n747_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n733_), .A2(new_n567_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n733_), .A2(KEYINPUT118), .A3(new_n567_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n765_), .A2(new_n768_), .A3(KEYINPUT58), .A4(new_n769_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n518_), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n752_), .A2(new_n764_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n762_), .B2(KEYINPUT57), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  INV_X1    g577(.A(new_n749_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n779_), .A2(new_n760_), .B1(new_n568_), .B2(new_n733_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT117), .B(new_n778_), .C1(new_n780_), .C2(new_n517_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n539_), .B1(new_n775_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n573_), .A2(new_n753_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT54), .B1(new_n658_), .B2(new_n784_), .ZN(new_n785_));
  OR4_X1    g584(.A1(KEYINPUT54), .A2(new_n518_), .A3(new_n539_), .A4(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n730_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n228_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT120), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n778_), .B1(new_n780_), .B2(new_n517_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n752_), .A2(new_n764_), .A3(new_n774_), .A4(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n539_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n787_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n730_), .A2(KEYINPUT59), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n788_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n796_), .B(KEYINPUT121), .C1(new_n788_), .C2(new_n797_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n753_), .A2(new_n266_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT122), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n790_), .B1(new_n802_), .B2(new_n804_), .ZN(G1340gat));
  OAI21_X1  g604(.A(G120gat), .B1(new_n798_), .B2(new_n575_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n262_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n788_), .B(new_n807_), .C1(KEYINPUT60), .C2(new_n262_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1341gat));
  NAND4_X1  g608(.A1(new_n800_), .A2(G127gat), .A3(new_n581_), .A4(new_n801_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n788_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n263_), .B1(new_n811_), .B2(new_n539_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1342gat));
  XNOR2_X1  g612(.A(KEYINPUT123), .B(G134gat), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n617_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n800_), .A2(new_n801_), .A3(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n264_), .B1(new_n811_), .B2(new_n580_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(KEYINPUT124), .A3(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1343gat));
  AOI211_X1 g621(.A(new_n284_), .B(new_n350_), .C1(new_n783_), .C2(new_n787_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n823_), .A2(new_n442_), .A3(new_n591_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n228_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n574_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n581_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  AOI21_X1  g630(.A(G162gat), .B1(new_n824_), .B2(new_n517_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n518_), .A2(G162gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT125), .Z(new_n834_));
  AOI21_X1  g633(.A(new_n832_), .B1(new_n824_), .B2(new_n834_), .ZN(G1347gat));
  NOR2_X1   g634(.A1(new_n591_), .A2(new_n442_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n284_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT126), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n794_), .A2(new_n350_), .A3(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G169gat), .B1(new_n839_), .B2(new_n753_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT62), .ZN(new_n841_));
  INV_X1    g640(.A(new_n839_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n228_), .A3(new_n355_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1348gat));
  NAND2_X1  g643(.A1(new_n783_), .A2(new_n787_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n845_), .A2(new_n350_), .A3(new_n838_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(G176gat), .A3(new_n574_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n235_), .B1(new_n839_), .B2(new_n573_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1349gat));
  AOI21_X1  g648(.A(G183gat), .B1(new_n846_), .B2(new_n581_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n364_), .A2(new_n247_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n839_), .A2(new_n539_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1350gat));
  OAI21_X1  g652(.A(G190gat), .B1(new_n839_), .B2(new_n617_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n517_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT127), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n839_), .B2(new_n856_), .ZN(G1351gat));
  NAND2_X1  g656(.A1(new_n823_), .A2(new_n836_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n753_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n575_), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g661(.A1(new_n858_), .A2(new_n539_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n863_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT63), .B(G211gat), .Z(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n863_), .B2(new_n865_), .ZN(G1354gat));
  NOR2_X1   g665(.A1(new_n858_), .A2(new_n580_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(G218gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n858_), .A2(new_n617_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(G218gat), .B2(new_n869_), .ZN(G1355gat));
endmodule


