//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_;
  NOR2_X1   g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(G57gat), .A2(G64gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT11), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  INV_X1    g007(.A(G71gat), .ZN(new_n209_));
  INV_X1    g008(.A(G78gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n206_), .A2(new_n208_), .A3(new_n212_), .A4(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n216_));
  OAI221_X1 g015(.A(KEYINPUT11), .B1(new_n207_), .B2(new_n202_), .C1(new_n211_), .C2(new_n213_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n216_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n220_), .B(new_n221_), .Z(new_n222_));
  XOR2_X1   g021(.A(G15gat), .B(G22gat), .Z(new_n223_));
  NAND2_X1  g022(.A1(G1gat), .A2(G8gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(KEYINPUT14), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT82), .ZN(new_n226_));
  XOR2_X1   g025(.A(G1gat), .B(G8gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n222_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT16), .B(G183gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(G211gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(G127gat), .B(G155gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT83), .Z(new_n237_));
  AND2_X1   g036(.A1(new_n233_), .A2(new_n234_), .ZN(new_n238_));
  OR3_X1    g037(.A1(new_n229_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241_));
  INV_X1    g040(.A(G99gat), .ZN(new_n242_));
  INV_X1    g041(.A(G106gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT6), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n244_), .A2(new_n247_), .A3(new_n248_), .A4(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(G85gat), .A2(G92gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G85gat), .A2(G92gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT67), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT8), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n250_), .A2(new_n259_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT64), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT9), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n251_), .A2(new_n263_), .A3(new_n265_), .A4(new_n252_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n263_), .A2(new_n252_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n247_), .A2(new_n248_), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT10), .B(G99gat), .Z(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n243_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n266_), .A2(new_n267_), .A3(KEYINPUT65), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n261_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT78), .B(G43gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G50gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G29gat), .B(G36gat), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n278_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT76), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT34), .ZN(new_n284_));
  OAI22_X1  g083(.A1(new_n276_), .A2(new_n281_), .B1(KEYINPUT35), .B2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n281_), .B(KEYINPUT15), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n285_), .B1(new_n287_), .B2(new_n276_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(KEYINPUT35), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT77), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n288_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT79), .B(G134gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G162gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT80), .B(KEYINPUT36), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT81), .Z(new_n298_));
  OR2_X1    g097(.A1(new_n291_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n295_), .B(KEYINPUT36), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n291_), .A2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT37), .Z(new_n303_));
  XNOR2_X1  g102(.A(G71gat), .B(G99gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G190gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT84), .B(G183gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT90), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT88), .Z(new_n316_));
  INV_X1    g115(.A(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT89), .B1(new_n318_), .B2(G169gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G169gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n317_), .B(new_n319_), .C1(new_n320_), .C2(KEYINPUT89), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n314_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT87), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(KEYINPUT24), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(new_n310_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n316_), .A2(KEYINPUT24), .A3(new_n324_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  OR3_X1    g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT25), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(KEYINPUT25), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n330_), .A2(new_n331_), .B1(KEYINPUT26), .B2(new_n311_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n312_), .A2(KEYINPUT25), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n311_), .A2(KEYINPUT26), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT86), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n327_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n322_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT91), .B(G113gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G120gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(G127gat), .B(G134gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n338_), .B(KEYINPUT30), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n344_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT31), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n346_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n307_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n346_), .A2(new_n348_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n350_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n346_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n306_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G141gat), .ZN(new_n363_));
  INV_X1    g162(.A(G148gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT92), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n365_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT2), .Z(new_n370_));
  OAI21_X1  g169(.A(new_n362_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n362_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n360_), .A2(KEYINPUT1), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(new_n369_), .A3(new_n365_), .A4(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT28), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n378_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G197gat), .ZN(new_n385_));
  INV_X1    g184(.A(G197gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(KEYINPUT21), .B2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n385_), .B(KEYINPUT94), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n387_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(KEYINPUT21), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT21), .A3(new_n383_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(new_n376_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n397_), .B(KEYINPUT93), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n394_), .B(new_n398_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT96), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n382_), .B1(new_n405_), .B2(KEYINPUT97), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n402_), .B(new_n404_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n359_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n354_), .A2(new_n358_), .A3(new_n408_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n344_), .B(new_n376_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT4), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OR3_X1    g215(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n376_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n414_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n415_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT0), .B(G57gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G85gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT105), .ZN(new_n426_));
  INV_X1    g225(.A(new_n424_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n418_), .A2(new_n419_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(KEYINPUT105), .A3(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(new_n338_), .B2(new_n394_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT19), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n316_), .B(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n320_), .A2(new_n317_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G183gat), .A2(G190gat), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n438_), .B(new_n439_), .C1(new_n310_), .C2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n324_), .A2(KEYINPUT24), .A3(new_n315_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT26), .B(G190gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT98), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT25), .B(G183gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n326_), .B(new_n442_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n433_), .B(new_n436_), .C1(new_n394_), .C2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n394_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n450_), .B(KEYINPUT20), .C1(new_n338_), .C2(new_n394_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n451_), .A2(KEYINPUT100), .A3(new_n435_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT100), .B1(new_n451_), .B2(new_n435_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G8gat), .B(G36gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  OR2_X1    g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n459_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT27), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n448_), .A2(KEYINPUT104), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT104), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n441_), .A2(new_n465_), .A3(new_n447_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n433_), .B1(new_n467_), .B2(new_n394_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n435_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n435_), .B2(new_n451_), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n459_), .B(KEYINPUT106), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n460_), .A2(new_n472_), .A3(KEYINPUT27), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n412_), .A2(new_n431_), .A3(new_n463_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n431_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n459_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT32), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n476_), .B(new_n480_), .C1(new_n454_), .C2(new_n479_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT102), .A2(KEYINPUT33), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n428_), .B(new_n482_), .Z(new_n483_));
  AND3_X1   g282(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n484_), .A2(KEYINPUT103), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n427_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(KEYINPUT103), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n460_), .A2(new_n483_), .A3(new_n461_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n481_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n359_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n409_), .A3(new_n491_), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n240_), .B(new_n303_), .C1(new_n475_), .C2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G230gat), .A2(G233gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n276_), .B2(new_n220_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT70), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n276_), .A2(new_n220_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n276_), .A2(KEYINPUT12), .A3(new_n220_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT70), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n495_), .C1(new_n276_), .C2(new_n220_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n498_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n276_), .A2(new_n220_), .ZN(new_n506_));
  OAI211_X1 g305(.A(G230gat), .B(G233gat), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT71), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G176gat), .B(G204gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT73), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n504_), .A2(new_n516_), .A3(new_n507_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n509_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT74), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n504_), .A2(new_n507_), .A3(new_n514_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT74), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n509_), .A2(new_n521_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT75), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n519_), .A2(KEYINPUT75), .A3(new_n520_), .A4(new_n522_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n494_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n494_), .A3(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n281_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n228_), .A2(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n226_), .A2(new_n227_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n226_), .A2(new_n227_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n281_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n533_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n228_), .A2(new_n534_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n540_), .B(new_n532_), .C1(new_n228_), .C2(new_n286_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G113gat), .B(G141gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(G169gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n386_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n539_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n531_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n493_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT107), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(G1gat), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n493_), .A2(new_n549_), .A3(KEYINPUT107), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n476_), .A4(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n555_), .A2(KEYINPUT108), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(KEYINPUT108), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT38), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n302_), .ZN(new_n560_));
  AOI211_X1 g359(.A(new_n240_), .B(new_n560_), .C1(new_n475_), .C2(new_n492_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n549_), .ZN(new_n562_));
  OAI21_X1  g361(.A(G1gat), .B1(new_n562_), .B2(new_n431_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT109), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n558_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n564_), .A3(new_n565_), .ZN(G1324gat));
  AND2_X1   g365(.A1(new_n552_), .A2(new_n554_), .ZN(new_n567_));
  INV_X1    g366(.A(G8gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n474_), .A2(new_n463_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n562_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(new_n569_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n572_), .A2(new_n573_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n570_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT40), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n570_), .B(KEYINPUT40), .C1(new_n575_), .C2(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(G1325gat));
  OAI21_X1  g380(.A(G15gat), .B1(new_n562_), .B2(new_n491_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT41), .Z(new_n583_));
  INV_X1    g382(.A(G15gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n567_), .A2(new_n584_), .A3(new_n359_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(G1326gat));
  INV_X1    g385(.A(G22gat), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n567_), .A2(new_n587_), .A3(new_n408_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G22gat), .B1(new_n562_), .B2(new_n409_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT110), .Z(new_n590_));
  AND2_X1   g389(.A1(new_n590_), .A2(KEYINPUT42), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(KEYINPUT42), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n588_), .B1(new_n591_), .B2(new_n592_), .ZN(G1327gat));
  AOI21_X1  g392(.A(new_n302_), .B1(new_n475_), .B2(new_n492_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n549_), .A2(new_n240_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n596_), .A2(G29gat), .A3(new_n431_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT44), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n302_), .B(KEYINPUT37), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n475_), .B2(new_n492_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT43), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n549_), .A2(new_n240_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n598_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT43), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n600_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n602_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(KEYINPUT44), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n476_), .A3(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n608_), .A2(KEYINPUT111), .A3(G29gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT111), .B1(new_n608_), .B2(G29gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n597_), .B1(new_n609_), .B2(new_n610_), .ZN(G1328gat));
  NAND2_X1  g410(.A1(new_n603_), .A2(new_n607_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n569_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G36gat), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(G36gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n595_), .A2(new_n615_), .A3(new_n569_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n614_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT46), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n614_), .A2(KEYINPUT46), .A3(new_n618_), .A4(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(G1329gat));
  NAND2_X1  g423(.A1(new_n359_), .A2(G43gat), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n596_), .A2(new_n491_), .ZN(new_n626_));
  OAI22_X1  g425(.A1(new_n612_), .A2(new_n625_), .B1(G43gat), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g427(.A(G50gat), .B1(new_n612_), .B2(new_n409_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n409_), .A2(G50gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT113), .Z(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n596_), .B2(new_n631_), .ZN(G1331gat));
  INV_X1    g431(.A(new_n548_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n530_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n561_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(G57gat), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n431_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT115), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n493_), .A2(new_n634_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n639_), .B2(new_n431_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT114), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n638_), .A2(new_n641_), .ZN(G1332gat));
  OAI21_X1  g441(.A(G64gat), .B1(new_n635_), .B2(new_n613_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT48), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n613_), .A2(G64gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n639_), .B2(new_n645_), .ZN(G1333gat));
  OAI21_X1  g445(.A(G71gat), .B1(new_n635_), .B2(new_n491_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT49), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n359_), .A2(new_n209_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n639_), .B2(new_n649_), .ZN(G1334gat));
  OAI21_X1  g449(.A(G78gat), .B1(new_n635_), .B2(new_n409_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT50), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n408_), .A2(new_n210_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n639_), .B2(new_n653_), .ZN(G1335gat));
  INV_X1    g453(.A(new_n240_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n530_), .A2(new_n633_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n594_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G85gat), .B1(new_n658_), .B2(new_n476_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n605_), .A2(G85gat), .A3(new_n656_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n476_), .ZN(G1336gat));
  NAND2_X1  g460(.A1(new_n605_), .A2(new_n656_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n569_), .A2(G92gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n657_), .A2(new_n613_), .ZN(new_n664_));
  OAI22_X1  g463(.A1(new_n662_), .A2(new_n663_), .B1(G92gat), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT116), .ZN(G1337gat));
  NAND3_X1  g465(.A1(new_n605_), .A2(new_n359_), .A3(new_n656_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G99gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT117), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT118), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT51), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n658_), .A2(new_n272_), .A3(new_n359_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .A4(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n668_), .A2(KEYINPUT117), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT117), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n667_), .B2(G99gat), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n670_), .B(new_n672_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT51), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n678_), .ZN(G1338gat));
  NAND3_X1  g478(.A1(new_n658_), .A2(new_n243_), .A3(new_n408_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n605_), .A2(new_n408_), .A3(new_n656_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT52), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G106gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G106gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g485(.A1(new_n569_), .A2(new_n431_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n410_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n546_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n532_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n540_), .B1(new_n228_), .B2(new_n286_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n692_), .B(new_n544_), .C1(new_n532_), .C2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT120), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n500_), .A2(new_n501_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n698_), .A2(KEYINPUT55), .A3(new_n497_), .A4(new_n503_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT55), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n504_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n500_), .A2(new_n501_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n506_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n699_), .B(new_n701_), .C1(new_n495_), .C2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n515_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n548_), .B1(new_n697_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT56), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT56), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n704_), .A2(KEYINPUT120), .A3(new_n708_), .A4(new_n515_), .ZN(new_n709_));
  AND4_X1   g508(.A1(new_n520_), .A2(new_n706_), .A3(new_n707_), .A4(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n302_), .B1(new_n696_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT57), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT57), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n302_), .C1(new_n696_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n695_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n704_), .A2(new_n708_), .A3(new_n515_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n716_), .A2(new_n520_), .A3(new_n707_), .A4(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT58), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n303_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n715_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT121), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n715_), .A2(KEYINPUT121), .A3(new_n720_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n240_), .A3(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n240_), .A2(new_n633_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n525_), .A2(new_n494_), .A3(new_n526_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n527_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT119), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT119), .B(new_n726_), .C1(new_n727_), .C2(new_n527_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n599_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT54), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT54), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n730_), .A2(new_n734_), .A3(new_n599_), .A4(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n690_), .B1(new_n725_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G113gat), .B1(new_n737_), .B2(new_n633_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n721_), .A2(new_n240_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT59), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n689_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n737_), .B2(new_n741_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n548_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n738_), .B1(new_n744_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g544(.A(G120gat), .B1(new_n743_), .B2(new_n530_), .ZN(new_n746_));
  INV_X1    g545(.A(G120gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n530_), .B2(KEYINPUT60), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n737_), .B(new_n748_), .C1(KEYINPUT60), .C2(new_n747_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1341gat));
  AOI21_X1  g549(.A(G127gat), .B1(new_n737_), .B2(new_n655_), .ZN(new_n751_));
  INV_X1    g550(.A(G127gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n743_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n753_), .B2(new_n655_), .ZN(G1342gat));
  NAND2_X1  g553(.A1(new_n737_), .A2(new_n560_), .ZN(new_n755_));
  INV_X1    g554(.A(G134gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT122), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT122), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n599_), .A2(new_n756_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n742_), .B(new_n761_), .C1(new_n737_), .C2(new_n741_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n758_), .A2(new_n760_), .A3(new_n762_), .ZN(G1343gat));
  AND2_X1   g562(.A1(new_n725_), .A2(new_n736_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n411_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n687_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G141gat), .B1(new_n766_), .B2(new_n548_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n764_), .A2(new_n411_), .A3(new_n688_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n363_), .A3(new_n633_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1344gat));
  OAI21_X1  g569(.A(G148gat), .B1(new_n766_), .B2(new_n530_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n364_), .A3(new_n531_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1345gat));
  NAND2_X1  g572(.A1(new_n725_), .A2(new_n736_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n411_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n774_), .A2(new_n655_), .A3(new_n775_), .A4(new_n687_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT61), .B(G155gat), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(G1346gat));
  NAND2_X1  g577(.A1(new_n768_), .A2(new_n560_), .ZN(new_n779_));
  INV_X1    g578(.A(G162gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n303_), .A2(G162gat), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT123), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n779_), .A2(new_n780_), .B1(new_n768_), .B2(new_n782_), .ZN(G1347gat));
  OAI211_X1 g582(.A(new_n431_), .B(new_n359_), .C1(new_n473_), .C2(new_n462_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT124), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n633_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n740_), .A2(new_n409_), .A3(new_n790_), .A4(new_n320_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT62), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(KEYINPUT125), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT125), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n788_), .A2(new_n794_), .A3(new_n633_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n408_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n740_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n792_), .B1(new_n797_), .B2(G169gat), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n733_), .A2(new_n735_), .B1(new_n240_), .B2(new_n721_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n794_), .B1(new_n788_), .B2(new_n633_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT125), .B(new_n548_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n409_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n792_), .B(G169gat), .C1(new_n799_), .C2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n791_), .B1(new_n798_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT126), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT126), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n791_), .C1(new_n798_), .C2(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(G1348gat));
  INV_X1    g608(.A(new_n788_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n799_), .A2(new_n408_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G176gat), .B1(new_n811_), .B2(new_n531_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n764_), .A2(new_n408_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n810_), .A2(new_n317_), .A3(new_n530_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(G1349gat));
  INV_X1    g614(.A(new_n811_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(new_n240_), .A3(new_n445_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n655_), .A3(new_n788_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n312_), .ZN(G1350gat));
  OAI21_X1  g618(.A(G190gat), .B1(new_n816_), .B2(new_n599_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n302_), .A2(new_n444_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n816_), .B2(new_n821_), .ZN(G1351gat));
  NAND2_X1  g621(.A1(new_n569_), .A2(new_n431_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n774_), .A2(new_n775_), .A3(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n548_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(KEYINPUT127), .A3(new_n386_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT127), .B(G197gat), .Z(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(new_n828_), .ZN(G1352gat));
  NOR2_X1   g628(.A1(new_n825_), .A2(new_n530_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(new_n384_), .ZN(G1353gat));
  XOR2_X1   g630(.A(KEYINPUT63), .B(G211gat), .Z(new_n832_));
  NAND4_X1  g631(.A1(new_n765_), .A2(new_n655_), .A3(new_n824_), .A4(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n825_), .B2(new_n240_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1354gat));
  INV_X1    g635(.A(G218gat), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n825_), .A2(new_n837_), .A3(new_n599_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n825_), .A2(new_n302_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n837_), .B2(new_n839_), .ZN(G1355gat));
endmodule


