//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT25), .B(G183gat), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n206_), .A2(G190gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(G190gat), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n212_), .A2(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n216_), .B(KEYINPUT23), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n213_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n211_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n215_), .A2(new_n220_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G197gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n227_), .A2(G204gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT88), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT21), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT88), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n227_), .B2(G204gat), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n229_), .B(new_n230_), .C1(new_n228_), .C2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G211gat), .B(G218gat), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G204gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G197gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n227_), .A2(G204gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT87), .B1(new_n239_), .B2(KEYINPUT21), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241_));
  AOI211_X1 g040(.A(new_n241_), .B(new_n230_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n233_), .B(new_n235_), .C1(new_n240_), .C2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n229_), .B1(new_n232_), .B2(new_n228_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(KEYINPUT21), .A3(new_n234_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT91), .B1(new_n243_), .B2(new_n245_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n226_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT20), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT98), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(KEYINPUT98), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n255_), .A2(KEYINPUT99), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT99), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n250_), .A2(new_n257_), .A3(new_n252_), .A4(new_n254_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT89), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n246_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n243_), .A2(KEYINPUT89), .A3(new_n245_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT26), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT80), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n266_), .A2(new_n267_), .B1(new_n205_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT80), .B1(new_n270_), .B2(G183gat), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n206_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT82), .B1(new_n272_), .B2(new_n207_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n218_), .A2(new_n275_), .A3(new_n219_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n212_), .A2(KEYINPUT24), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT83), .B1(new_n221_), .B2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n279_), .A3(new_n214_), .ZN(new_n280_));
  AOI21_X1  g079(.A(G183gat), .B1(new_n263_), .B2(new_n264_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n225_), .B1(new_n218_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n262_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n258_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n204_), .B1(new_n256_), .B2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n260_), .A2(new_n280_), .A3(new_n261_), .A4(new_n282_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT20), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT96), .ZN(new_n289_));
  INV_X1    g088(.A(new_n204_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n246_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n226_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT96), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n287_), .A2(new_n294_), .A3(KEYINPUT20), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n289_), .A2(new_n290_), .A3(new_n293_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n286_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G92gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT18), .B(G64gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n202_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n226_), .A2(new_n291_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n290_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n289_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n204_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT101), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n287_), .A2(new_n294_), .A3(KEYINPUT20), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n294_), .B1(new_n287_), .B2(KEYINPUT20), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n313_), .A2(new_n314_), .A3(new_n292_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n305_), .B1(new_n315_), .B2(new_n290_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n302_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n202_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n303_), .A2(KEYINPUT101), .A3(new_n309_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n312_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT2), .ZN(new_n325_));
  INV_X1    g124(.A(G141gat), .ZN(new_n326_));
  INV_X1    g125(.A(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT86), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n326_), .B(new_n327_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT85), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(KEYINPUT1), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n328_), .B(new_n324_), .C1(new_n337_), .C2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n323_), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n262_), .A2(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G78gat), .B(G106gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT92), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n248_), .A2(new_n249_), .A3(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n345_), .B(new_n348_), .C1(new_n351_), .C2(new_n322_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT93), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n345_), .B1(new_n351_), .B2(new_n322_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n347_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n353_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n343_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(G50gat), .B1(new_n343_), .B2(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT28), .B(G22gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n362_), .A3(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n352_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n355_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT94), .B1(new_n370_), .B2(new_n346_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n352_), .A2(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  INV_X1    g172(.A(new_n346_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n355_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n367_), .A2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G127gat), .B(G134gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XOR2_X1   g179(.A(G113gat), .B(G120gat), .Z(new_n381_));
  XNOR2_X1  g180(.A(G127gat), .B(G134gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n380_), .A2(new_n383_), .A3(KEYINPUT84), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT84), .B1(new_n380_), .B2(new_n383_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n386_), .B(KEYINPUT30), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(new_n283_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT31), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n388_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n391_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n386_), .A2(new_n343_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n340_), .A2(new_n380_), .A3(new_n383_), .A4(new_n342_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT4), .B1(new_n386_), .B2(new_n343_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n396_), .A3(new_n400_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n403_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n395_), .A2(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n321_), .A2(new_n377_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n301_), .A2(KEYINPUT32), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n297_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n412_), .B1(new_n308_), .B2(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n403_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n396_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n399_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n408_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT97), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT33), .A4(new_n409_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n425_), .A2(new_n426_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n317_), .A2(new_n429_), .A3(new_n309_), .A4(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n419_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT100), .B1(new_n432_), .B2(new_n377_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n377_), .B1(new_n419_), .B2(new_n431_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT100), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n312_), .A2(new_n377_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n412_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n433_), .B(new_n436_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n395_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT66), .ZN(new_n442_));
  NAND3_X1  g241(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(KEYINPUT66), .A3(new_n443_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G92gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n452_), .A2(G92gat), .ZN(new_n455_));
  OAI21_X1  g254(.A(G85gat), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G85gat), .B(G92gat), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT9), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT10), .B(G99gat), .Z(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n451_), .A2(new_n456_), .A3(new_n458_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT68), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT67), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n444_), .A2(new_n445_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n460_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n464_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n457_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT8), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n457_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n465_), .A2(new_n466_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n451_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n463_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n477_), .B1(new_n474_), .B2(new_n457_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n483_), .A2(KEYINPUT68), .A3(new_n480_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n462_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n488_), .A2(new_n489_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(KEYINPUT12), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G230gat), .A2(G233gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n495_), .B(KEYINPUT64), .Z(new_n496_));
  OAI21_X1  g295(.A(new_n462_), .B1(new_n483_), .B2(new_n480_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n493_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n494_), .A2(new_n496_), .A3(new_n498_), .A4(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n499_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G204gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT5), .B(G176gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n510_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(new_n505_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(KEYINPUT13), .A3(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n520_));
  XNOR2_X1  g319(.A(G29gat), .B(G36gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G29gat), .B(G36gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n522_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n519_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n525_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n522_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(KEYINPUT15), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G15gat), .ZN(new_n535_));
  INV_X1    g334(.A(G22gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G15gat), .A2(G22gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G1gat), .A2(G8gat), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n537_), .A2(new_n538_), .B1(KEYINPUT14), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(G1gat), .A2(G8gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT76), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n539_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n542_), .B2(new_n539_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n541_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n529_), .A2(new_n534_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n549_), .B(new_n547_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G169gat), .B(G197gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n558_), .A3(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n518_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n441_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT36), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT72), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(KEYINPUT72), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n529_), .A2(new_n534_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n476_), .A2(new_n463_), .A3(new_n481_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT68), .B1(new_n483_), .B2(new_n480_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n581_), .B1(new_n584_), .B2(new_n462_), .ZN(new_n585_));
  OAI221_X1 g384(.A(new_n462_), .B1(new_n527_), .B2(new_n528_), .C1(new_n483_), .C2(new_n480_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n576_), .A2(new_n577_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n579_), .B(new_n580_), .C1(new_n585_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n581_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n485_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n588_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n591_), .A2(KEYINPUT72), .A3(new_n578_), .A4(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n589_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n573_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT74), .B(new_n573_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n589_), .A2(new_n593_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n572_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .A4(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n492_), .B(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n550_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT78), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n613_), .B(new_n619_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n611_), .A2(KEYINPUT17), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT79), .Z(new_n623_));
  NAND4_X1  g422(.A1(new_n599_), .A2(new_n603_), .A3(new_n606_), .A4(new_n600_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n589_), .A2(new_n593_), .A3(new_n573_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n606_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n602_), .B1(new_n626_), .B2(KEYINPUT37), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n607_), .A2(new_n623_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n569_), .A2(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n630_), .A2(G1gat), .A3(new_n412_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT38), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n599_), .A2(new_n606_), .A3(new_n600_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT102), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n599_), .A2(new_n635_), .A3(new_n606_), .A4(new_n600_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n569_), .A2(new_n622_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n638_), .B2(new_n412_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n631_), .A2(KEYINPUT38), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n632_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT103), .ZN(G1324gat));
  INV_X1    g441(.A(new_n630_), .ZN(new_n643_));
  INV_X1    g442(.A(G8gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n321_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n569_), .A2(new_n622_), .A3(new_n637_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n321_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n648_), .B2(G8gat), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT39), .B(new_n644_), .C1(new_n647_), .C2(new_n321_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n645_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1325gat));
  NAND3_X1  g452(.A1(new_n643_), .A2(new_n535_), .A3(new_n395_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n647_), .A2(new_n395_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(G15gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n655_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n535_), .B(new_n658_), .C1(new_n647_), .C2(new_n395_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(KEYINPUT41), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT41), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n654_), .B1(new_n661_), .B2(new_n662_), .ZN(G1326gat));
  XNOR2_X1  g462(.A(new_n377_), .B(KEYINPUT106), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G22gat), .B1(new_n638_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n643_), .A2(new_n536_), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n637_), .A2(new_n623_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n434_), .B(KEYINPUT100), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n303_), .A2(KEYINPUT101), .A3(new_n309_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT101), .B1(new_n303_), .B2(new_n309_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n412_), .A3(new_n377_), .A4(new_n319_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n395_), .B1(new_n671_), .B2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n567_), .B(new_n670_), .C1(new_n676_), .C2(new_n414_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n439_), .A2(new_n440_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n414_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n682_), .A2(KEYINPUT107), .A3(new_n567_), .A4(new_n670_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n679_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n438_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n624_), .A2(new_n627_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n624_), .A2(KEYINPUT75), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n441_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT43), .B(new_n691_), .C1(new_n676_), .C2(new_n414_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n623_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n690_), .A2(new_n567_), .A3(new_n692_), .A4(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(KEYINPUT44), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n697_), .A2(G29gat), .A3(new_n438_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(KEYINPUT44), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n685_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n679_), .A2(new_n683_), .A3(new_n702_), .A4(new_n321_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n321_), .B1(new_n694_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G36gat), .B1(new_n696_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n684_), .A2(new_n710_), .A3(new_n702_), .A4(new_n321_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(KEYINPUT45), .A3(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n709_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n706_), .A2(new_n713_), .A3(new_n709_), .A4(KEYINPUT46), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n694_), .B2(new_n707_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n699_), .A2(new_n395_), .A3(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n684_), .A2(new_n395_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(G43gat), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n684_), .B2(new_n664_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n699_), .A2(G50gat), .A3(new_n377_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n697_), .ZN(G1331gat));
  INV_X1    g526(.A(new_n566_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n518_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n441_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n629_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT109), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n438_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n637_), .A3(new_n623_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT110), .B1(new_n438_), .B2(G57gat), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(G57gat), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n734_), .A2(KEYINPUT110), .A3(new_n735_), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n733_), .A2(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(new_n321_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G64gat), .B1(new_n734_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT48), .ZN(new_n742_));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n743_), .A3(new_n321_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n734_), .B2(new_n440_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n732_), .A2(new_n748_), .A3(new_n395_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1334gat));
  NOR2_X1   g549(.A1(new_n665_), .A2(G78gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT112), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n732_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G78gat), .B1(new_n734_), .B2(new_n665_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT111), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(KEYINPUT111), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n758_), .B2(new_n759_), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n729_), .A2(new_n728_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n682_), .A2(new_n670_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT113), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n682_), .A2(new_n764_), .A3(new_n670_), .A4(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n438_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n690_), .A2(new_n693_), .A3(new_n692_), .A4(new_n761_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n438_), .A2(G85gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n766_), .B2(new_n321_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n455_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n740_), .B1(new_n773_), .B2(new_n453_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n769_), .B2(new_n774_), .ZN(G1337gat));
  OAI21_X1  g574(.A(G99gat), .B1(new_n768_), .B2(new_n440_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n766_), .A2(new_n459_), .A3(new_n395_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779_));
  INV_X1    g578(.A(new_n459_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(new_n395_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT115), .B(new_n776_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT51), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n777_), .A2(KEYINPUT114), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n779_), .A3(new_n395_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n787_), .A2(KEYINPUT115), .A3(new_n788_), .A4(new_n776_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n784_), .A2(new_n789_), .ZN(G1338gat));
  INV_X1    g589(.A(new_n377_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G106gat), .B1(new_n768_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT52), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(G106gat), .C1(new_n768_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n766_), .A2(new_n460_), .A3(new_n377_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT53), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n800_), .A3(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n634_), .A2(new_n636_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n494_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n504_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT55), .A3(new_n502_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n502_), .A2(KEYINPUT55), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n510_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n807_), .A2(new_n808_), .A3(new_n811_), .A4(new_n510_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n810_), .A2(new_n728_), .A3(new_n513_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n551_), .A2(new_n557_), .A3(new_n553_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n556_), .A2(new_n552_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n562_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n565_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n565_), .A2(new_n817_), .A3(KEYINPUT116), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n814_), .B1(new_n514_), .B2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n502_), .A2(new_n505_), .A3(new_n512_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n512_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n814_), .B(new_n822_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n813_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n803_), .B1(new_n804_), .B2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n810_), .A2(new_n513_), .A3(new_n812_), .A4(new_n822_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n812_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n805_), .B2(new_n504_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n512_), .B1(new_n836_), .B2(new_n502_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n811_), .B1(new_n837_), .B2(new_n808_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n513_), .A4(new_n822_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n833_), .B(new_n840_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n830_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT119), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n813_), .A2(new_n828_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n637_), .A2(new_n844_), .A3(KEYINPUT57), .A4(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n845_), .A2(KEYINPUT57), .A3(new_n634_), .A4(new_n636_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT118), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n830_), .A2(new_n841_), .A3(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n843_), .A2(new_n849_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n693_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n629_), .A2(new_n854_), .A3(new_n566_), .A4(new_n729_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n607_), .A2(new_n566_), .A3(new_n623_), .A4(new_n628_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n856_), .B2(new_n518_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n321_), .A2(new_n412_), .A3(new_n377_), .A4(new_n440_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n842_), .B1(new_n848_), .B2(new_n846_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n858_), .B1(new_n863_), .B2(new_n622_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT59), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n728_), .B2(G113gat), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n728_), .B(new_n872_), .C1(new_n867_), .C2(new_n869_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(G1340gat));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n729_), .B2(G120gat), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n872_), .B(new_n876_), .C1(new_n875_), .C2(G120gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G120gat), .B1(new_n867_), .B2(new_n729_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n872_), .B2(new_n623_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n867_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n622_), .A2(G127gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n872_), .B2(new_n804_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT122), .B(G134gat), .Z(new_n887_));
  NOR2_X1   g686(.A1(new_n689_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n883_), .B2(new_n888_), .ZN(G1343gat));
  AND2_X1   g688(.A1(new_n864_), .A2(new_n438_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n437_), .A2(new_n395_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n566_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n326_), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n729_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n327_), .ZN(G1345gat));
  NOR2_X1   g695(.A1(new_n892_), .A2(new_n693_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT61), .B(G155gat), .Z(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  INV_X1    g698(.A(G162gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n892_), .A2(new_n900_), .A3(new_n689_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n890_), .A2(new_n804_), .A3(new_n891_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n900_), .B2(new_n902_), .ZN(G1347gat));
  AND2_X1   g702(.A1(new_n728_), .A2(new_n224_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n740_), .A2(new_n413_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n665_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n859_), .B2(new_n908_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n855_), .A2(new_n857_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n852_), .B2(new_n693_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n911_), .A2(KEYINPUT124), .A3(new_n907_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n904_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n842_), .A2(KEYINPUT119), .B1(new_n848_), .B2(new_n846_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n623_), .B1(new_n914_), .B2(new_n851_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n728_), .B(new_n908_), .C1(new_n915_), .C2(new_n910_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G169gat), .ZN(new_n917_));
  OR2_X1    g716(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n918_));
  NAND2_X1  g717(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n916_), .A2(KEYINPUT123), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n913_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT125), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n913_), .A2(new_n920_), .A3(new_n924_), .A4(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1348gat));
  OR2_X1    g725(.A1(new_n909_), .A2(new_n912_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n518_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n864_), .A2(new_n791_), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n740_), .A2(new_n211_), .A3(new_n729_), .A4(new_n413_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n928_), .A2(new_n211_), .B1(new_n929_), .B2(new_n930_), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n623_), .A3(new_n906_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT126), .ZN(new_n933_));
  INV_X1    g732(.A(G183gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n622_), .A2(new_n205_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n934_), .B1(new_n927_), .B2(new_n935_), .ZN(G1350gat));
  NAND2_X1  g735(.A1(new_n927_), .A2(new_n691_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G190gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n207_), .A2(new_n208_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n927_), .A2(new_n939_), .A3(new_n804_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1351gat));
  AND2_X1   g740(.A1(new_n864_), .A2(new_n440_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n740_), .A2(new_n438_), .A3(new_n791_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n566_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n227_), .ZN(G1352gat));
  INV_X1    g745(.A(new_n944_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n518_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n236_), .A2(KEYINPUT127), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1353gat));
  AOI211_X1 g749(.A(KEYINPUT63), .B(G211gat), .C1(new_n947_), .C2(new_n622_), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT63), .B(G211gat), .Z(new_n952_));
  AND3_X1   g751(.A1(new_n947_), .A2(new_n622_), .A3(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n944_), .A2(new_n955_), .A3(new_n689_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n947_), .A2(new_n804_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n955_), .B2(new_n957_), .ZN(G1355gat));
endmodule


