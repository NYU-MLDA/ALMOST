//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G232gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT34), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n205_), .B2(KEYINPUT35), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G36gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G29gat), .ZN(new_n210_));
  INV_X1    g009(.A(G29gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G36gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n208_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n211_), .A2(G36gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n209_), .A2(G29gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT74), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(new_n207_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT15), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n235_), .A3(KEYINPUT67), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n242_));
  NOR2_X1   g041(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n232_), .B2(new_n235_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT8), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n241_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n249_));
  OAI22_X1  g048(.A1(new_n246_), .A2(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(new_n240_), .ZN(new_n252_));
  OR2_X1    g051(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n251_), .A2(new_n239_), .A3(new_n240_), .A4(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n252_), .A2(new_n257_), .A3(new_n259_), .A4(new_n235_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n250_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n206_), .B1(new_n226_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n205_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT35), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n232_), .A2(new_n235_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(new_n236_), .A3(new_n245_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n232_), .A2(new_n235_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT8), .B1(new_n272_), .B2(new_n241_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n267_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n222_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n262_), .A2(new_n266_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n206_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n223_), .A2(new_n225_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n274_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n261_), .A2(new_n222_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n265_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G190gat), .B(G218gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT36), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(new_n282_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n285_), .B(KEYINPUT36), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n289_), .B2(KEYINPUT76), .ZN(new_n290_));
  INV_X1    g089(.A(new_n288_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n266_), .B1(new_n262_), .B2(new_n276_), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n280_), .A2(new_n281_), .A3(new_n265_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n202_), .B(KEYINPUT37), .C1(new_n290_), .C2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n298_), .A2(KEYINPUT37), .A3(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n295_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n289_), .A2(KEYINPUT76), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n287_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n202_), .B1(new_n303_), .B2(KEYINPUT37), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G15gat), .B(G22gat), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G8gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G71gat), .B(G78gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G57gat), .B(G64gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(KEYINPUT11), .B2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n316_), .A2(KEYINPUT11), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(KEYINPUT11), .ZN(new_n320_));
  INV_X1    g119(.A(new_n315_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n314_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G155gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G183gat), .B(G211gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT17), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n329_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n333_), .B1(new_n331_), .B2(new_n323_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n305_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT79), .ZN(new_n337_));
  XOR2_X1   g136(.A(KEYINPUT89), .B(G204gat), .Z(new_n338_));
  INV_X1    g137(.A(KEYINPUT90), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(G197gat), .ZN(new_n340_));
  INV_X1    g139(.A(G204gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n341_), .B2(G197gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT89), .B(G204gat), .ZN(new_n343_));
  INV_X1    g142(.A(G197gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n340_), .A2(KEYINPUT92), .A3(new_n345_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G211gat), .B(G218gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n338_), .A2(G197gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n344_), .A2(G204gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT21), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n340_), .A2(new_n345_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n360_), .A3(new_n351_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(KEYINPUT87), .A3(new_n366_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(KEYINPUT2), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G141gat), .A2(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT3), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n373_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n371_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n377_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n366_), .B1(new_n364_), .B2(KEYINPUT1), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n385_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT88), .B1(new_n384_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n369_), .A2(new_n370_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n383_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n375_), .A2(new_n378_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n390_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n362_), .B(new_n363_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n384_), .A2(new_n391_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n353_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n358_), .A2(new_n360_), .A3(new_n351_), .ZN(new_n406_));
  OAI22_X1  g205(.A1(new_n404_), .A2(new_n402_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n363_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(KEYINPUT94), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n401_), .A2(new_n402_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT28), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT28), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n401_), .A2(new_n418_), .A3(new_n402_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G22gat), .B(G50gat), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n423_));
  AOI211_X1 g222(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n392_), .C2(new_n400_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n420_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n403_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n415_), .A2(new_n422_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n410_), .A2(new_n411_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n403_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n403_), .A2(new_n409_), .A3(KEYINPUT93), .A4(new_n412_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G127gat), .B(G134gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G113gat), .B(G120gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT23), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(G183gat), .B2(G190gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT83), .Z(new_n445_));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n446_));
  INV_X1    g245(.A(G169gat), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT22), .ZN(new_n448_));
  INV_X1    g247(.A(G176gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT22), .B1(new_n446_), .B2(new_n447_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n445_), .A3(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G169gat), .A2(G176gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n445_), .A2(KEYINPUT24), .A3(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT25), .B(G183gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT26), .B(G190gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n442_), .B(new_n459_), .C1(new_n455_), .C2(KEYINPUT24), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n452_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT30), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464_));
  INV_X1    g263(.A(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G227gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(G15gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n466_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n463_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT31), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n461_), .A2(new_n462_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(new_n462_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n470_), .A3(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n472_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n440_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n476_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n470_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT31), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n472_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n439_), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n436_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n484_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(new_n427_), .C1(new_n430_), .C2(new_n435_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n392_), .A2(new_n400_), .A3(new_n440_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n404_), .A2(new_n439_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n439_), .A2(KEYINPUT4), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n392_), .A2(new_n400_), .A3(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n497_), .A2(new_n494_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(KEYINPUT4), .A3(new_n491_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT95), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n502_), .A3(new_n499_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n495_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G57gat), .B(G85gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT97), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G1gat), .B(G29gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT98), .B1(new_n504_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n495_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n503_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n502_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT98), .ZN(new_n516_));
  INV_X1    g315(.A(new_n510_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n512_), .B(new_n510_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n511_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n455_), .A2(KEYINPUT24), .A3(new_n444_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n453_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n521_), .A2(new_n442_), .A3(new_n459_), .A4(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT22), .B(G169gat), .Z(new_n525_));
  OAI211_X1 g324(.A(new_n443_), .B(new_n445_), .C1(G176gat), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT20), .B(new_n528_), .C1(new_n362_), .C2(new_n461_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G226gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT19), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n362_), .A2(new_n461_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n355_), .A2(new_n361_), .A3(new_n526_), .A4(new_n524_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n533_), .A2(KEYINPUT20), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G8gat), .B(G36gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT18), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G64gat), .B(G92gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n529_), .A2(new_n534_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n540_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n533_), .A2(KEYINPUT20), .A3(new_n535_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n544_), .B(new_n545_), .C1(new_n534_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n541_), .A2(new_n542_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT27), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n532_), .A2(new_n536_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT27), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n541_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n489_), .A2(new_n520_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n511_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n544_), .B1(new_n546_), .B2(new_n534_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n540_), .A2(KEYINPUT32), .ZN(new_n559_));
  MUX2_X1   g358(.A(new_n558_), .B(new_n551_), .S(new_n559_), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n519_), .A2(KEYINPUT33), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n504_), .A2(new_n562_), .A3(new_n510_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n499_), .A2(new_n493_), .A3(new_n497_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(new_n517_), .C1(new_n493_), .C2(new_n492_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n552_), .A2(new_n541_), .A3(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n557_), .A2(new_n560_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n436_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n485_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n556_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n312_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT81), .B1(new_n573_), .B2(new_n275_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT81), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n312_), .A2(new_n222_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n275_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT80), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n574_), .A2(KEYINPUT80), .A3(new_n578_), .A4(new_n576_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n578_), .B1(new_n279_), .B2(new_n573_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n581_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n586_), .A3(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n322_), .B1(new_n250_), .B2(new_n260_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT12), .B1(new_n595_), .B2(KEYINPUT69), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n250_), .A2(new_n260_), .A3(new_n322_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT64), .Z(new_n600_));
  INV_X1    g399(.A(KEYINPUT69), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n601_), .B(new_n602_), .C1(new_n274_), .C2(new_n322_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n596_), .A2(new_n598_), .A3(new_n600_), .A4(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G176gat), .B(G204gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT71), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n600_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n597_), .B2(new_n595_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT72), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n604_), .A2(new_n612_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n610_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(KEYINPUT72), .A3(new_n613_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n621_));
  OR2_X1    g420(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n622_));
  NAND2_X1  g421(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n617_), .A2(new_n619_), .A3(new_n622_), .A4(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n572_), .A2(new_n594_), .A3(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n337_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n307_), .A3(new_n557_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT101), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n557_), .A2(new_n560_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n564_), .A2(new_n567_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n486_), .A2(new_n488_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n635_), .A2(new_n570_), .B1(new_n636_), .B2(new_n520_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n298_), .A2(new_n289_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT100), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n594_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n625_), .A2(new_n334_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n520_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n632_), .B(new_n645_), .C1(new_n630_), .C2(new_n629_), .ZN(G1324gat));
  INV_X1    g445(.A(new_n555_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n647_), .A3(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n628_), .A2(new_n308_), .A3(new_n647_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n644_), .B2(new_n487_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n628_), .A2(new_n468_), .A3(new_n485_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n644_), .B2(new_n436_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n628_), .A2(new_n666_), .A3(new_n569_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1327gat));
  NOR2_X1   g467(.A1(new_n639_), .A2(new_n335_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n627_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n557_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n300_), .A2(KEYINPUT104), .A3(new_n304_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT43), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n673_), .B1(new_n637_), .B2(new_n305_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n300_), .A2(new_n304_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(KEYINPUT43), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n572_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n621_), .A2(new_n334_), .A3(new_n594_), .A4(new_n624_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT103), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT44), .B1(new_n678_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n683_), .B(new_n680_), .C1(new_n674_), .C2(new_n677_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n520_), .A2(new_n211_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n671_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n670_), .A2(new_n209_), .A3(new_n647_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n685_), .B2(new_n647_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n572_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n676_), .B1(new_n572_), .B2(new_n675_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n681_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n683_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT44), .B(new_n681_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n695_), .A2(KEYINPUT105), .A3(new_n647_), .A4(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n690_), .B1(new_n691_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n690_), .B(KEYINPUT46), .C1(new_n691_), .C2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1329gat));
  NAND2_X1  g502(.A1(new_n695_), .A2(new_n696_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G43gat), .B1(new_n704_), .B2(new_n487_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n670_), .A2(new_n465_), .A3(new_n485_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1330gat));
  OAI21_X1  g508(.A(G50gat), .B1(new_n704_), .B2(new_n436_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n436_), .A2(G50gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT107), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n670_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1331gat));
  AOI21_X1  g513(.A(new_n594_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n641_), .A2(new_n335_), .A3(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(G57gat), .A3(new_n557_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n637_), .B2(new_n594_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n572_), .A2(new_n719_), .A3(new_n642_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n718_), .A2(new_n625_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n337_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(new_n520_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n723_), .B2(G57gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT109), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n716_), .A2(new_n647_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G64gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n555_), .A2(G64gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n722_), .B2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n716_), .B2(new_n485_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n485_), .A2(new_n732_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n722_), .B2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n716_), .B2(new_n569_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT50), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n569_), .A2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n722_), .B2(new_n740_), .ZN(G1335gat));
  NAND4_X1  g540(.A1(new_n718_), .A2(new_n625_), .A3(new_n669_), .A4(new_n720_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n237_), .A3(new_n557_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n715_), .A2(new_n334_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT111), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n678_), .A2(KEYINPUT112), .A3(new_n746_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n520_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n744_), .B1(new_n751_), .B2(new_n237_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT113), .ZN(G1336gat));
  NAND3_X1  g552(.A1(new_n743_), .A2(new_n238_), .A3(new_n647_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n555_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n238_), .ZN(G1337gat));
  OR2_X1    g555(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n757_));
  NAND2_X1  g556(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n485_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n742_), .A2(KEYINPUT114), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT114), .B1(new_n742_), .B2(new_n759_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n749_), .A2(new_n750_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n227_), .B1(new_n764_), .B2(new_n485_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n757_), .B(new_n758_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n485_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G99gat), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n762_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n766_), .A2(new_n769_), .ZN(G1338gat));
  NAND4_X1  g569(.A1(new_n743_), .A2(new_n254_), .A3(new_n256_), .A4(new_n569_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n678_), .A2(new_n569_), .A3(new_n746_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n772_), .A2(new_n773_), .A3(G106gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n772_), .B2(G106gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g576(.A(new_n582_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n590_), .B1(new_n585_), .B2(new_n581_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n587_), .B2(new_n591_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n617_), .A2(new_n781_), .A3(new_n619_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n604_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n322_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT69), .B1(new_n261_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n597_), .B1(new_n786_), .B2(new_n602_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n787_), .A2(KEYINPUT55), .A3(new_n600_), .A4(new_n596_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n603_), .A2(new_n598_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n261_), .A2(new_n785_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n602_), .B1(new_n790_), .B2(new_n601_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n611_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n784_), .A2(new_n788_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n616_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n615_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n592_), .A2(new_n593_), .B1(new_n799_), .B2(new_n610_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n793_), .A2(new_n795_), .A3(new_n616_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n782_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n639_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(new_n639_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n616_), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n809_), .A2(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(KEYINPUT119), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n781_), .A2(new_n613_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT58), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n812_), .B1(new_n809_), .B2(KEYINPUT119), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n817_), .B(KEYINPUT56), .C1(new_n793_), .C2(new_n616_), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT58), .B(new_n814_), .C1(new_n816_), .C2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n675_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n807_), .A2(new_n808_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n814_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n675_), .A3(new_n819_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n826_), .B(new_n827_), .C1(new_n808_), .C2(new_n807_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n335_), .B1(new_n822_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n642_), .A2(new_n335_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT116), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n626_), .A2(new_n831_), .A3(new_n305_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n829_), .A2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n647_), .A2(new_n520_), .A3(new_n486_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n594_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(G113gat), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n821_), .A2(new_n334_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n835_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n838_), .B1(new_n829_), .B2(new_n836_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(KEYINPUT59), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n594_), .A2(new_n847_), .A3(G113gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n847_), .B2(G113gat), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n839_), .A2(new_n840_), .B1(new_n846_), .B2(new_n849_), .ZN(G1340gat));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n846_), .B2(new_n625_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n625_), .A2(new_n854_), .A3(new_n852_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n845_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n853_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n857_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n626_), .B(new_n844_), .C1(new_n845_), .C2(KEYINPUT59), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n859_), .B(KEYINPUT122), .C1(new_n860_), .C2(new_n852_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(G1341gat));
  AND2_X1   g661(.A1(new_n846_), .A2(new_n335_), .ZN(new_n863_));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n335_), .A2(new_n864_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n863_), .A2(new_n864_), .B1(new_n845_), .B2(new_n865_), .ZN(G1342gat));
  AND2_X1   g665(.A1(new_n846_), .A2(new_n675_), .ZN(new_n867_));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n640_), .A2(new_n868_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n867_), .A2(new_n868_), .B1(new_n845_), .B2(new_n869_), .ZN(G1343gat));
  INV_X1    g669(.A(new_n488_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n647_), .A2(new_n520_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n837_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n642_), .ZN(new_n874_));
  INV_X1    g673(.A(G141gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1344gat));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n626_), .ZN(new_n877_));
  INV_X1    g676(.A(G148gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n873_), .A2(new_n334_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n873_), .B2(new_n305_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n639_), .A2(G162gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n873_), .B2(new_n884_), .ZN(G1347gat));
  NAND2_X1  g684(.A1(new_n835_), .A2(new_n843_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n555_), .A2(new_n557_), .A3(new_n486_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G169gat), .B1(new_n888_), .B2(new_n642_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n890_));
  OR2_X1    g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n890_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n642_), .A2(new_n525_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT124), .Z(new_n894_));
  OAI211_X1 g693(.A(new_n891_), .B(new_n892_), .C1(new_n888_), .C2(new_n894_), .ZN(G1348gat));
  INV_X1    g694(.A(new_n888_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n896_), .B2(new_n625_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n887_), .A2(G176gat), .A3(new_n625_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n837_), .B2(new_n898_), .ZN(G1349gat));
  NOR2_X1   g698(.A1(new_n888_), .A2(new_n334_), .ZN(new_n900_));
  MUX2_X1   g699(.A(G183gat), .B(new_n457_), .S(new_n900_), .Z(G1350gat));
  NAND3_X1  g700(.A1(new_n896_), .A2(new_n458_), .A3(new_n640_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n896_), .A2(new_n675_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n903_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(KEYINPUT125), .B1(new_n903_), .B2(G190gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1351gat));
  NOR2_X1   g705(.A1(new_n555_), .A2(new_n557_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n871_), .B(new_n907_), .C1(new_n829_), .C2(new_n836_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n642_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n344_), .ZN(G1352gat));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n626_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n338_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n341_), .B2(new_n911_), .ZN(G1353gat));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NOR4_X1   g714(.A1(new_n908_), .A2(new_n334_), .A3(new_n914_), .A4(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n908_), .B2(new_n334_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n918_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n916_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  OAI21_X1  g720(.A(G218gat), .B1(new_n908_), .B2(new_n305_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n639_), .A2(G218gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n908_), .B2(new_n923_), .ZN(G1355gat));
endmodule


