//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_;
  XOR2_X1   g000(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT20), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT82), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n213_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT90), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(new_n213_), .C1(new_n216_), .C2(new_n218_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  MUX2_X1   g024(.A(new_n223_), .B(new_n224_), .S(new_n225_), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n214_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G169gat), .ZN(new_n230_));
  INV_X1    g029(.A(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n217_), .B(KEYINPUT83), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT91), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT91), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(KEYINPUT23), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n223_), .A2(new_n225_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(KEYINPUT85), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n237_), .A2(KEYINPUT85), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n235_), .B(new_n236_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n229_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G197gat), .B(G204gat), .Z(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT21), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(KEYINPUT21), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n210_), .B1(new_n244_), .B2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n232_), .B(new_n233_), .C1(new_n226_), .C2(new_n242_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n254_), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT25), .B1(new_n254_), .B2(G183gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n211_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OAI221_X1 g056(.A(new_n257_), .B1(KEYINPUT24), .B2(new_n215_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n215_), .A2(KEYINPUT24), .A3(new_n233_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(new_n251_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n209_), .B1(new_n252_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n210_), .B1(new_n260_), .B2(new_n251_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n229_), .A2(new_n249_), .A3(new_n250_), .A4(new_n243_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n263_), .A2(new_n209_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266_));
  NOR3_X1   g065(.A1(new_n262_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n209_), .A3(new_n264_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(KEYINPUT92), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n206_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n244_), .A2(new_n251_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n261_), .A2(new_n271_), .A3(KEYINPUT20), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n268_), .B(KEYINPUT92), .C1(new_n272_), .C2(new_n209_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n206_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n269_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n276_), .A3(KEYINPUT94), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n267_), .A2(new_n269_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT94), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n274_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n278_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n209_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n272_), .B2(new_n209_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n270_), .B(KEYINPUT27), .C1(new_n206_), .C2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT2), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(KEYINPUT2), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT3), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(KEYINPUT3), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n301_), .B2(new_n297_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n292_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n289_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT29), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n251_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G78gat), .B(G106gat), .Z(new_n313_));
  AOI22_X1  g112(.A1(new_n307_), .A2(new_n251_), .B1(new_n310_), .B2(new_n309_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n312_), .B(new_n313_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT89), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n312_), .B1(new_n314_), .B2(new_n311_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n306_), .A2(KEYINPUT29), .ZN(new_n320_));
  XOR2_X1   g119(.A(G22gat), .B(G50gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n320_), .B(new_n323_), .ZN(new_n324_));
  AND4_X1   g123(.A1(new_n315_), .A2(new_n316_), .A3(new_n319_), .A4(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n316_), .A2(new_n324_), .B1(new_n319_), .B2(new_n315_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n306_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n300_), .A2(new_n330_), .A3(new_n305_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT95), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT95), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n332_), .A2(new_n340_), .A3(KEYINPUT4), .A4(new_n333_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n332_), .ZN(new_n342_));
  XOR2_X1   g141(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n343_));
  AOI22_X1  g142(.A1(new_n339_), .A2(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n335_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n337_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n347_));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G57gat), .B(G85gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(new_n345_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n336_), .A3(new_n351_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G71gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n330_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT30), .B(G99gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G15gat), .B(G43gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT31), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n260_), .B(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n361_), .B(new_n364_), .Z(new_n365_));
  NOR2_X1   g164(.A1(new_n355_), .A2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n286_), .A2(new_n327_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT33), .B1(new_n346_), .B2(new_n351_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n344_), .A2(new_n335_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n351_), .B1(new_n334_), .B2(new_n345_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n354_), .B2(new_n372_), .ZN(new_n373_));
  AOI211_X1 g172(.A(new_n368_), .B(new_n373_), .C1(new_n277_), .C2(new_n281_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n352_), .A2(new_n354_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n273_), .A2(new_n275_), .B1(KEYINPUT32), .B2(new_n206_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n284_), .A2(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n375_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n327_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n355_), .A2(new_n327_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n282_), .A3(new_n285_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT98), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT98), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n381_), .A2(new_n282_), .A3(new_n384_), .A4(new_n285_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n367_), .B1(new_n386_), .B2(new_n365_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT5), .B(G176gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G204gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G120gat), .B(G148gat), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(KEYINPUT68), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT69), .Z(new_n394_));
  NAND2_X1  g193(.A1(G230gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT64), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT6), .ZN(new_n401_));
  AND2_X1   g200(.A1(G99gat), .A2(G106gat), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n402_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n397_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G99gat), .A2(G106gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n400_), .A2(KEYINPUT6), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n398_), .A2(KEYINPUT64), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(KEYINPUT65), .A3(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G85gat), .B(G92gat), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT8), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n415_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n417_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT8), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n405_), .A2(new_n411_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT9), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n418_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(G85gat), .A3(G92gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT10), .B(G99gat), .Z(new_n430_));
  INV_X1    g229(.A(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .A4(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT66), .B(G71gat), .ZN(new_n434_));
  INV_X1    g233(.A(G78gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G57gat), .B(G64gat), .Z(new_n437_));
  INV_X1    g236(.A(KEYINPUT11), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n434_), .B(G78gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n424_), .A2(new_n433_), .A3(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n442_), .A2(new_n444_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n416_), .A2(new_n419_), .B1(new_n422_), .B2(KEYINPUT8), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n405_), .A2(new_n411_), .A3(new_n429_), .A4(new_n432_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(new_n427_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n447_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n451_), .A3(KEYINPUT12), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n424_), .A2(new_n433_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n447_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n396_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n395_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT67), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n457_), .A2(KEYINPUT67), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n394_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n394_), .B1(new_n459_), .B2(new_n458_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT13), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT13), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G43gat), .B(G50gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n466_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT15), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n474_), .A2(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n472_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT79), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT77), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n472_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n485_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n481_), .A2(KEYINPUT77), .A3(new_n472_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n490_), .A2(KEYINPUT78), .A3(new_n491_), .A4(new_n492_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n487_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G113gat), .B(G141gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n487_), .A2(new_n495_), .A3(new_n496_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(KEYINPUT80), .A3(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n465_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n387_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n453_), .A2(new_n474_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n513_), .B(new_n518_), .C1(new_n472_), .C2(new_n453_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n516_), .A2(new_n517_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT71), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(KEYINPUT36), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT71), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n526_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT37), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n527_), .A2(new_n529_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(KEYINPUT72), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n481_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n447_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT73), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G127gat), .B(G155gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT16), .B(G183gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(KEYINPUT73), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n544_), .A2(KEYINPUT17), .A3(new_n548_), .A4(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT74), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT74), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n543_), .B(KEYINPUT75), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n548_), .B(KEYINPUT17), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT76), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n540_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n512_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n476_), .A3(new_n355_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT38), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT99), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n510_), .A2(new_n557_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(new_n534_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n386_), .A2(new_n365_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n367_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n566_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n476_), .B1(new_n574_), .B2(new_n355_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n564_), .A2(new_n576_), .ZN(G1324gat));
  OAI21_X1  g376(.A(G8gat), .B1(new_n573_), .B2(new_n286_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT101), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT101), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(G8gat), .C1(new_n573_), .C2(new_n286_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(KEYINPUT39), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n286_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n560_), .A2(new_n477_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(KEYINPUT101), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(G1325gat));
  OAI21_X1  g388(.A(G15gat), .B1(new_n573_), .B2(new_n365_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G15gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n365_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n560_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n595_), .ZN(G1326gat));
  INV_X1    g395(.A(G22gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n327_), .B(KEYINPUT103), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n560_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT42), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n574_), .A2(new_n599_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n602_), .B2(G22gat), .ZN(new_n603_));
  AOI211_X1 g402(.A(KEYINPUT42), .B(new_n597_), .C1(new_n574_), .C2(new_n599_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT104), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  NOR2_X1   g408(.A1(new_n557_), .A2(new_n538_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n512_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G29gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n355_), .A2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT106), .Z(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT44), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n571_), .A2(new_n617_), .A3(new_n540_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n540_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT43), .B1(new_n387_), .B2(new_n619_), .ZN(new_n620_));
  AOI211_X1 g419(.A(new_n511_), .B(new_n557_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n616_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n620_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n510_), .A3(new_n558_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n375_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n615_), .B1(new_n627_), .B2(new_n612_), .ZN(G1328gat));
  INV_X1    g427(.A(G36gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n611_), .A2(new_n629_), .A3(new_n583_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(new_n632_));
  AOI21_X1  g431(.A(new_n286_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(new_n629_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n632_), .B(new_n635_), .C1(new_n633_), .C2(new_n629_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1329gat));
  INV_X1    g438(.A(G43gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n611_), .A2(new_n640_), .A3(new_n594_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n365_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n640_), .ZN(new_n643_));
  XOR2_X1   g442(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n644_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n646_), .B(new_n641_), .C1(new_n642_), .C2(new_n640_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1330gat));
  INV_X1    g447(.A(G50gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n611_), .A2(new_n649_), .A3(new_n599_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n327_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(new_n649_), .ZN(G1331gat));
  INV_X1    g451(.A(new_n465_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n387_), .A2(new_n508_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n559_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n355_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n654_), .A2(new_n538_), .A3(new_n557_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(new_n355_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n659_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g459(.A(G64gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n658_), .B2(new_n583_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT48), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(new_n661_), .A3(new_n583_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1333gat));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n356_), .A3(new_n594_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n594_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G71gat), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n668_), .A2(KEYINPUT111), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(KEYINPUT111), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n666_), .B1(new_n672_), .B2(new_n673_), .ZN(G1334gat));
  AOI21_X1  g473(.A(new_n435_), .B1(new_n658_), .B2(new_n599_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT50), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n656_), .A2(new_n435_), .A3(new_n599_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1335gat));
  NOR2_X1   g477(.A1(new_n653_), .A2(new_n508_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n558_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT112), .Z(new_n682_));
  OAI21_X1  g481(.A(G85gat), .B1(new_n682_), .B2(new_n375_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n654_), .A2(new_n610_), .ZN(new_n684_));
  INV_X1    g483(.A(G85gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n355_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(G1336gat));
  OAI21_X1  g486(.A(G92gat), .B1(new_n682_), .B2(new_n286_), .ZN(new_n688_));
  INV_X1    g487(.A(G92gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n684_), .A2(new_n689_), .A3(new_n583_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1337gat));
  NAND2_X1  g490(.A1(new_n681_), .A2(new_n594_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G99gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n430_), .A3(new_n594_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT113), .A3(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1338gat));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n327_), .B(new_n680_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(KEYINPUT115), .A3(new_n431_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT115), .ZN(new_n701_));
  INV_X1    g500(.A(new_n327_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n680_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n624_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n704_), .B2(G106gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n700_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT115), .B1(new_n699_), .B2(new_n431_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n701_), .A3(G106gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(KEYINPUT52), .A3(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n684_), .A2(new_n431_), .A3(new_n702_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n706_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n706_), .A2(new_n709_), .A3(new_n710_), .A4(new_n712_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1339gat));
  NAND3_X1  g515(.A1(new_n458_), .A2(new_n392_), .A3(new_n459_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n508_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT118), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n452_), .A2(new_n396_), .A3(new_n455_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT55), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n456_), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT55), .B(new_n396_), .C1(new_n452_), .C2(new_n455_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n452_), .A2(new_n455_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n395_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(KEYINPUT55), .A3(new_n720_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n723_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(KEYINPUT118), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n724_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT56), .B1(new_n730_), .B2(new_n391_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT56), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n732_), .B(new_n392_), .C1(new_n724_), .C2(new_n729_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n718_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT119), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n490_), .A2(new_n486_), .A3(new_n492_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n484_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n736_), .B(new_n500_), .C1(new_n737_), .C2(new_n486_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(new_n503_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n462_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT119), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n741_), .B(new_n718_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n735_), .A2(new_n740_), .A3(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(KEYINPUT57), .A3(new_n538_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT120), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n538_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT57), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n731_), .A2(new_n733_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n739_), .A3(new_n717_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n749_), .A2(KEYINPUT58), .A3(new_n739_), .A4(new_n717_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n540_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT120), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n743_), .A2(new_n755_), .A3(KEYINPUT57), .A4(new_n538_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n745_), .A2(new_n748_), .A3(new_n754_), .A4(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n558_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  AND4_X1   g559(.A1(new_n509_), .A2(new_n536_), .A3(new_n539_), .A4(new_n557_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n653_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n536_), .A2(new_n539_), .A3(new_n509_), .A4(new_n557_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n763_), .A2(new_n465_), .A3(KEYINPUT117), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n760_), .A3(new_n653_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT117), .B1(new_n763_), .B2(new_n465_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(KEYINPUT54), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n758_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n583_), .A2(new_n702_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n355_), .A3(new_n594_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(KEYINPUT121), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT121), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n769_), .B1(new_n757_), .B2(new_n558_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n773_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G113gat), .B1(new_n779_), .B2(new_n508_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n771_), .A2(new_n781_), .A3(new_n774_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT59), .B1(new_n777_), .B2(new_n773_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(new_n509_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n780_), .B1(G113gat), .B2(new_n785_), .ZN(G1340gat));
  INV_X1    g585(.A(G120gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n653_), .B2(KEYINPUT60), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n779_), .B(new_n788_), .C1(KEYINPUT60), .C2(new_n787_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G120gat), .B1(new_n784_), .B2(new_n653_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1341gat));
  NAND4_X1  g590(.A1(new_n782_), .A2(new_n783_), .A3(G127gat), .A4(new_n557_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n558_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G127gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT122), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT122), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n792_), .C1(new_n793_), .C2(G127gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1342gat));
  AOI21_X1  g597(.A(G134gat), .B1(new_n779_), .B2(new_n534_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n784_), .A2(new_n619_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(G134gat), .B2(new_n800_), .ZN(G1343gat));
  NOR3_X1   g600(.A1(new_n777_), .A2(new_n375_), .A3(new_n594_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n583_), .A2(new_n327_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n508_), .A3(new_n803_), .ZN(new_n804_));
  XOR2_X1   g603(.A(KEYINPUT123), .B(G141gat), .Z(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1344gat));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n465_), .A3(new_n803_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT124), .B(G148gat), .Z(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1345gat));
  NAND3_X1  g608(.A1(new_n802_), .A2(new_n557_), .A3(new_n803_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT61), .B(G155gat), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1346gat));
  AND4_X1   g611(.A1(G162gat), .A2(new_n802_), .A3(new_n540_), .A4(new_n803_), .ZN(new_n813_));
  INV_X1    g612(.A(G162gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n802_), .A2(new_n534_), .A3(new_n803_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(G1347gat));
  INV_X1    g615(.A(KEYINPUT62), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n777_), .A2(new_n599_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n583_), .A2(new_n366_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n509_), .ZN(new_n822_));
  INV_X1    g621(.A(G169gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n817_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n230_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT62), .B(G169gat), .C1(new_n821_), .C2(new_n509_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(G1348gat));
  INV_X1    g626(.A(new_n821_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G176gat), .B1(new_n828_), .B2(new_n465_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n777_), .A2(new_n231_), .A3(new_n653_), .A4(new_n702_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n820_), .B2(new_n830_), .ZN(G1349gat));
  NAND4_X1  g630(.A1(new_n771_), .A2(new_n327_), .A3(new_n557_), .A4(new_n820_), .ZN(new_n832_));
  INV_X1    g631(.A(G183gat), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n819_), .A2(new_n212_), .A3(new_n558_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n832_), .A2(new_n833_), .B1(new_n818_), .B2(new_n834_), .ZN(G1350gat));
  OAI21_X1  g634(.A(G190gat), .B1(new_n821_), .B2(new_n619_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n534_), .A2(new_n211_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n821_), .B2(new_n837_), .ZN(G1351gat));
  INV_X1    g637(.A(new_n381_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n777_), .A2(new_n286_), .A3(new_n594_), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n508_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n465_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g643(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n771_), .A2(new_n583_), .A3(new_n365_), .A4(new_n381_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n558_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n845_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n845_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n840_), .A2(new_n850_), .A3(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1354gat));
  AOI21_X1  g656(.A(G218gat), .B1(new_n840_), .B2(new_n534_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n540_), .A2(G218gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT127), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n858_), .B1(new_n840_), .B2(new_n860_), .ZN(G1355gat));
endmodule


