//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  NOR2_X1   g000(.A1(G85gat), .A2(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n202_), .B1(new_n205_), .B2(KEYINPUT9), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G85gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n207_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n204_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n215_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n206_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  AOI211_X1 g021(.A(new_n218_), .B(new_n220_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI22_X1  g029(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n227_), .A2(new_n230_), .A3(new_n219_), .A4(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n220_), .A2(new_n218_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(KEYINPUT67), .A3(new_n231_), .A4(new_n227_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n205_), .A2(KEYINPUT8), .A3(new_n202_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n205_), .A2(new_n202_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(KEYINPUT68), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT8), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n232_), .B2(new_n239_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n238_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G29gat), .B(G36gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G43gat), .B(G50gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n224_), .A2(new_n243_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT34), .Z(new_n249_));
  INV_X1    g048(.A(KEYINPUT35), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT75), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n232_), .A2(new_n239_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT8), .A3(new_n240_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n256_), .A2(new_n238_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G29gat), .B(G36gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(new_n245_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT15), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT15), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n246_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n247_), .B(new_n252_), .C1(new_n257_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT77), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT76), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n224_), .A2(new_n243_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT76), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n247_), .A4(new_n252_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n249_), .A2(new_n250_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n266_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OAI221_X1 g071(.A(KEYINPUT76), .B1(new_n250_), .B2(new_n249_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT78), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n274_), .A2(KEYINPUT78), .A3(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT79), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n272_), .A2(new_n285_), .A3(new_n273_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n277_), .B(KEYINPUT36), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n285_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n284_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n291_), .A2(KEYINPUT80), .A3(new_n286_), .A4(new_n287_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n283_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT37), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n272_), .A2(new_n273_), .A3(new_n287_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT37), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT81), .B(G1gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT82), .B(G8gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT14), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G8gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n305_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(new_n303_), .B2(KEYINPUT14), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G57gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(G64gat), .ZN(new_n315_));
  INV_X1    g114(.A(G64gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(G57gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT11), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n315_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G71gat), .B(G78gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT69), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(G57gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(G64gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT11), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n321_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n319_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n320_), .A2(new_n322_), .A3(KEYINPUT69), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n327_), .B1(new_n326_), .B2(new_n321_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n319_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n313_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G231gat), .A2(G233gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT83), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n335_), .B(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G127gat), .B(G155gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(G183gat), .B(G211gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT17), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT85), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n343_), .A2(KEYINPUT17), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n300_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT1), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT97), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n353_), .B1(new_n356_), .B2(KEYINPUT1), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT96), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n357_), .A2(new_n358_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n355_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT95), .ZN(new_n364_));
  NOR2_X1   g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT98), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n365_), .B(KEYINPUT3), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n368_), .B(new_n369_), .C1(KEYINPUT2), .C2(new_n364_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n356_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n353_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT99), .Z(new_n373_));
  AOI22_X1  g172(.A1(new_n362_), .A2(new_n366_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(new_n370_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n366_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n378_), .B(new_n376_), .C1(new_n361_), .C2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT28), .ZN(new_n381_));
  XOR2_X1   g180(.A(G22gat), .B(G50gat), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n377_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n352_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n381_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n382_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n377_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n352_), .A2(KEYINPUT101), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n378_), .B1(new_n361_), .B2(new_n379_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT29), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G197gat), .B(G204gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(G211gat), .B(G218gat), .Z(new_n395_));
  INV_X1    g194(.A(KEYINPUT21), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n396_), .B2(new_n395_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n395_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n394_), .A3(KEYINPUT21), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n393_), .A2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(G228gat), .A2(G233gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n398_), .A2(KEYINPUT100), .A3(new_n400_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT100), .B1(new_n398_), .B2(new_n400_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(new_n403_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n393_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n404_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n386_), .A2(new_n391_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n386_), .B2(new_n391_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G113gat), .B(G120gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT90), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(G169gat), .B2(G176gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT24), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT23), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT91), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n429_), .A3(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G169gat), .A2(G176gat), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n419_), .A2(KEYINPUT24), .A3(new_n421_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT89), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G190gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(KEYINPUT26), .Z(new_n435_));
  INV_X1    g234(.A(KEYINPUT25), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT88), .A3(G183gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT25), .B(G183gat), .Z(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n438_), .B2(KEYINPUT88), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .A4(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n426_), .B1(G183gat), .B2(G190gat), .ZN(new_n442_));
  INV_X1    g241(.A(G176gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT22), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(KEYINPUT92), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G169gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n445_), .A2(G169gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT30), .B1(new_n441_), .B2(new_n448_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT93), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G43gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n451_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G43gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458_));
  INV_X1    g257(.A(G15gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n453_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n462_));
  OAI22_X1  g261(.A1(new_n449_), .A2(new_n450_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n441_), .A2(new_n448_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n461_), .A2(new_n462_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n441_), .A2(KEYINPUT30), .A3(new_n448_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT31), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n463_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n463_), .B2(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n417_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT31), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n463_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n416_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n473_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n413_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n386_), .A2(new_n391_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n410_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n386_), .A2(new_n391_), .A3(new_n410_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n473_), .A2(new_n477_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n481_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT27), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n448_), .B(new_n441_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n492_));
  XOR2_X1   g291(.A(KEYINPUT22), .B(G169gat), .Z(new_n493_));
  OAI211_X1 g292(.A(new_n442_), .B(new_n431_), .C1(G176gat), .C2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT25), .B(G183gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT26), .B(G190gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n424_), .A2(new_n426_), .A3(new_n432_), .A4(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n401_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT102), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT102), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n494_), .A2(new_n498_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n503_), .B2(new_n401_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n492_), .B(KEYINPUT20), .C1(new_n501_), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G226gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT19), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n507_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n464_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n510_), .B(new_n511_), .C1(new_n407_), .C2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G8gat), .B(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT18), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G64gat), .B(G92gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  AND3_X1   g316(.A1(new_n508_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n491_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n508_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n505_), .A2(new_n511_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n507_), .B(new_n510_), .C1(new_n407_), .C2(new_n512_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n521_), .B(KEYINPUT27), .C1(new_n524_), .C2(new_n517_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G225gat), .A2(G233gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT103), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n374_), .A2(new_n530_), .A3(new_n417_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n378_), .B(new_n530_), .C1(new_n361_), .C2(new_n379_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n416_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n374_), .A2(KEYINPUT4), .A3(new_n416_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n528_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G29gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT0), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n314_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(new_n203_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n533_), .A3(new_n527_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n536_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT104), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT104), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n542_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n526_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n517_), .A2(KEYINPUT32), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n524_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n508_), .A2(new_n513_), .A3(new_n550_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n551_), .B(new_n552_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n536_), .A2(new_n541_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n540_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(KEYINPUT33), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n531_), .A2(new_n533_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT4), .ZN(new_n558_));
  INV_X1    g357(.A(new_n535_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n528_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n527_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n540_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n519_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n556_), .A2(new_n562_), .A3(new_n521_), .A4(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n544_), .A2(KEYINPUT33), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n553_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n487_), .A2(KEYINPUT94), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n473_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n413_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n490_), .A2(new_n549_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n224_), .A2(new_n334_), .A3(new_n243_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n334_), .B1(new_n243_), .B2(new_n224_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(KEYINPUT70), .ZN(new_n575_));
  INV_X1    g374(.A(new_n334_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n267_), .A2(KEYINPUT70), .A3(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT12), .B1(new_n574_), .B2(KEYINPUT71), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n580_), .B(new_n581_), .C1(new_n257_), .C2(new_n334_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n579_), .A2(new_n571_), .A3(new_n573_), .A4(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G176gat), .B(G204gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT73), .ZN(new_n585_));
  XOR2_X1   g384(.A(G120gat), .B(G148gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n578_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT74), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n578_), .A2(new_n583_), .A3(new_n592_), .A4(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n578_), .A2(new_n583_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n589_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n594_), .A2(KEYINPUT13), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT13), .B1(new_n594_), .B2(new_n597_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n309_), .A2(KEYINPUT86), .A3(new_n259_), .A4(new_n312_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT86), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n313_), .B2(new_n246_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n259_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n602_), .B(new_n603_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n312_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n311_), .A2(new_n307_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n246_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n309_), .A2(new_n260_), .A3(new_n262_), .A4(new_n312_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n601_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT87), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT87), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n610_), .A2(new_n611_), .A3(new_n614_), .A4(new_n601_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G169gat), .B(G197gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n616_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n600_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n570_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n351_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n545_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n548_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OR3_X1    g428(.A1(new_n625_), .A2(new_n301_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n631_), .A2(KEYINPUT38), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT106), .ZN(new_n633_));
  INV_X1    g432(.A(new_n293_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n570_), .A2(new_n634_), .A3(new_n350_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT105), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n623_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n600_), .A2(KEYINPUT105), .A3(new_n622_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n628_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n631_), .A2(KEYINPUT38), .B1(new_n642_), .B2(G1gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n633_), .A2(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(new_n526_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G8gat), .B1(new_n640_), .B2(new_n645_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n646_), .A2(KEYINPUT107), .A3(KEYINPUT39), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT107), .B1(new_n646_), .B2(KEYINPUT39), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(KEYINPUT39), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n625_), .A2(new_n302_), .A3(new_n645_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n650_), .A2(KEYINPUT40), .A3(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  NAND2_X1  g455(.A1(new_n567_), .A2(new_n568_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n459_), .B1(new_n641_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n459_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n661_), .B(new_n662_), .C1(new_n625_), .C2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n640_), .B2(new_n486_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n486_), .A2(G22gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT108), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n625_), .B2(new_n668_), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n293_), .A2(new_n349_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n624_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n628_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n349_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n298_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n570_), .B2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(KEYINPUT43), .C1(new_n570_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n490_), .A2(new_n549_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n566_), .A2(new_n569_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n300_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n679_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT44), .B(new_n674_), .C1(new_n677_), .C2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n679_), .A3(new_n684_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n689_), .B2(new_n674_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT110), .A3(new_n628_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT110), .B1(new_n691_), .B2(new_n628_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n673_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  INV_X1    g495(.A(G36gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n691_), .B2(new_n526_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n671_), .A2(new_n697_), .A3(new_n526_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n687_), .A2(new_n690_), .A3(new_n645_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n702_), .B(KEYINPUT46), .C1(new_n697_), .C2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1329gat));
  NAND3_X1  g504(.A1(new_n671_), .A2(new_n456_), .A3(new_n658_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n687_), .A2(new_n690_), .A3(new_n487_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n456_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT47), .B(new_n706_), .C1(new_n707_), .C2(new_n456_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n671_), .B2(new_n413_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n413_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n691_), .B2(new_n714_), .ZN(G1331gat));
  NOR3_X1   g514(.A1(new_n570_), .A2(new_n622_), .A3(new_n600_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n351_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n628_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n720_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n293_), .A3(new_n349_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n723_), .A2(new_n314_), .A3(new_n629_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n721_), .A2(new_n722_), .A3(new_n724_), .ZN(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n723_), .B2(new_n645_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n727_));
  OR2_X1    g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n718_), .A2(new_n316_), .A3(new_n526_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n723_), .B2(new_n657_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT49), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n657_), .A2(G71gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n717_), .B2(new_n734_), .ZN(G1334gat));
  OAI21_X1  g534(.A(G78gat), .B1(new_n723_), .B2(new_n486_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT50), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n486_), .A2(G78gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n717_), .B2(new_n738_), .ZN(G1335gat));
  NAND2_X1  g538(.A1(new_n716_), .A2(new_n670_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n203_), .B1(new_n740_), .B2(new_n629_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT113), .Z(new_n742_));
  INV_X1    g541(.A(new_n600_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n350_), .A3(new_n621_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT114), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n689_), .A2(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n628_), .A2(new_n211_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n746_), .B2(new_n747_), .ZN(G1336gat));
  OAI21_X1  g547(.A(new_n204_), .B1(new_n740_), .B2(new_n645_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT115), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n645_), .A2(new_n204_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n746_), .B2(new_n751_), .ZN(G1337gat));
  INV_X1    g551(.A(new_n740_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n753_), .A2(new_n221_), .A3(new_n488_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n746_), .A2(new_n658_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G99gat), .ZN(new_n756_));
  XOR2_X1   g555(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1338gat));
  NAND3_X1  g557(.A1(new_n753_), .A2(new_n222_), .A3(new_n413_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n689_), .A2(new_n413_), .A3(new_n745_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G106gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G106gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g564(.A1(new_n675_), .A2(new_n349_), .A3(new_n621_), .A4(new_n600_), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n621_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n583_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n573_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT71), .B1(new_n267_), .B2(new_n576_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n581_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n776_), .A2(KEYINPUT55), .A3(new_n571_), .A4(new_n579_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n582_), .A2(new_n573_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n267_), .A2(new_n576_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n581_), .B1(new_n779_), .B2(new_n580_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n572_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(new_n777_), .A3(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n596_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n771_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n594_), .A2(new_n597_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n616_), .A2(new_n619_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n610_), .A2(new_n611_), .A3(new_n602_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n619_), .B(new_n788_), .C1(new_n789_), .C2(new_n602_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n787_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n785_), .A2(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(KEYINPUT118), .A3(new_n293_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT118), .B1(new_n793_), .B2(new_n293_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n770_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n594_), .A2(new_n791_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n782_), .A2(new_n596_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n594_), .A2(KEYINPUT120), .A3(new_n791_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n799_), .A2(new_n804_), .A3(new_n810_), .A4(new_n805_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n288_), .A2(new_n289_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n812_), .A2(KEYINPUT80), .B1(new_n281_), .B2(new_n282_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT37), .B1(new_n813_), .B2(new_n290_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n809_), .B(new_n811_), .C1(new_n814_), .C2(new_n298_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n793_), .A2(KEYINPUT57), .A3(new_n293_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n796_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n769_), .B1(new_n817_), .B2(new_n349_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n629_), .A2(new_n526_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n413_), .A2(new_n487_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(new_n819_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n816_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n815_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n796_), .A2(KEYINPUT119), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n300_), .A2(KEYINPUT122), .A3(new_n809_), .A4(new_n811_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n770_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .A4(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n768_), .B1(new_n832_), .B2(new_n350_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n822_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n824_), .B(new_n622_), .C1(new_n834_), .C2(new_n819_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G113gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n828_), .A2(new_n831_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n815_), .A2(new_n826_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n829_), .A3(new_n816_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n350_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n769_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n823_), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n842_), .A2(G113gat), .A3(new_n621_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n836_), .A2(new_n843_), .ZN(G1340gat));
  OAI211_X1 g643(.A(new_n824_), .B(new_n743_), .C1(new_n834_), .C2(new_n819_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT123), .B(G120gat), .Z(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n743_), .A2(new_n849_), .A3(new_n846_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n849_), .B2(new_n846_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n834_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n852_), .ZN(G1341gat));
  OAI211_X1 g652(.A(new_n824_), .B(new_n349_), .C1(new_n834_), .C2(new_n819_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G127gat), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n842_), .A2(G127gat), .A3(new_n350_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1342gat));
  NOR3_X1   g656(.A1(new_n833_), .A2(new_n293_), .A3(new_n822_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT124), .B1(new_n858_), .B2(G134gat), .ZN(new_n859_));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n675_), .A2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n824_), .B(new_n861_), .C1(new_n834_), .C2(new_n819_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n841_), .A2(new_n634_), .A3(new_n823_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n860_), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n859_), .A2(new_n862_), .A3(new_n865_), .ZN(G1343gat));
  INV_X1    g665(.A(new_n481_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n820_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n840_), .B2(new_n769_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n622_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n743_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT125), .B(G148gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1345gat));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n869_), .B2(new_n349_), .ZN(new_n877_));
  NOR4_X1   g676(.A1(new_n833_), .A2(KEYINPUT126), .A3(new_n350_), .A4(new_n868_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n868_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n793_), .A2(new_n293_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n793_), .A2(KEYINPUT118), .A3(new_n293_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n830_), .B1(new_n885_), .B2(new_n770_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n831_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n838_), .A2(new_n829_), .A3(new_n816_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n349_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n349_), .B(new_n880_), .C1(new_n890_), .C2(new_n768_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT126), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n869_), .A2(new_n876_), .A3(new_n349_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n875_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n879_), .A2(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(new_n869_), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n897_), .A2(G162gat), .A3(new_n293_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G162gat), .B1(new_n897_), .B2(new_n675_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1347gat));
  NAND3_X1  g699(.A1(new_n629_), .A2(new_n658_), .A3(new_n526_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT127), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n413_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n818_), .A2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G169gat), .B1(new_n904_), .B2(new_n621_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI211_X1 g706(.A(KEYINPUT62), .B(G169gat), .C1(new_n904_), .C2(new_n621_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n904_), .A2(new_n621_), .A3(new_n493_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1348gat));
  NOR2_X1   g709(.A1(new_n833_), .A2(new_n413_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n902_), .A2(new_n443_), .A3(new_n600_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n818_), .A2(new_n743_), .A3(new_n903_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n911_), .A2(new_n912_), .B1(new_n913_), .B2(new_n443_), .ZN(G1349gat));
  NOR3_X1   g713(.A1(new_n904_), .A2(new_n350_), .A3(new_n495_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n902_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n349_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(G183gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n904_), .B2(new_n675_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n634_), .A2(new_n496_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n904_), .B2(new_n921_), .ZN(G1351gat));
  NOR3_X1   g721(.A1(new_n628_), .A2(new_n481_), .A3(new_n645_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n841_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925_), .B2(new_n622_), .ZN(new_n926_));
  INV_X1    g725(.A(G197gat), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n924_), .A2(new_n927_), .A3(new_n621_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1352gat));
  OR3_X1    g728(.A1(new_n924_), .A2(G204gat), .A3(new_n600_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G204gat), .B1(new_n924_), .B2(new_n600_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1353gat));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n349_), .A2(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n925_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n936_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n924_), .A2(new_n933_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1354gat));
  OR3_X1    g739(.A1(new_n924_), .A2(G218gat), .A3(new_n293_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G218gat), .B1(new_n924_), .B2(new_n675_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(G1355gat));
endmodule


